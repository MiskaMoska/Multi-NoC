`timescale 1ns/1ns
`include "uvm_macros.svh"

import uvm_pkg::*;
`include "param.vh"
`include "cibd_if.sv"
`include "cibd_transaction.sv"
`include "cibd_driver.sv"
`include "cibd_monitor.sv"
`include "cibd_sequencer.sv"
`include "cibd_agent.sv"
`include "nop_model.sv"
`include "nop_scoreboard.sv"
`include "nop_env.sv"
`include "nop_base_test.sv"
`include "nop_sequence.sv"
`include "nop_case0.sv"

module top_tb;
reg clk_d;
reg clk_p;
reg rstn;

cibd_if i_if[75](clk_d,rstn);
cibd_if o_if[75](clk_d,rstn);

NoP dut(
    .CDCLK                           (clk_d),
    .CPCLK                           (clk_p),
    .CDRESETn                        (rstn),
    .CDIDATA_X0_Y0_D0                (i_if[0].data),
    .CDIVALID_X0_Y0_D0               (i_if[0].valid),
    .CDIREADY_X0_Y0_D0               (i_if[0].ready),
    .CDODATA_X0_Y0_D0                (o_if[0].data),
    .CDOVALID_X0_Y0_D0               (o_if[0].valid),
    .CDOREADY_X0_Y0_D0               (o_if[0].ready),

    .CDIDATA_X0_Y1_D0                (i_if[1].data),
    .CDIVALID_X0_Y1_D0               (i_if[1].valid),
    .CDIREADY_X0_Y1_D0               (i_if[1].ready),
    .CDODATA_X0_Y1_D0                (o_if[1].data),
    .CDOVALID_X0_Y1_D0               (o_if[1].valid),
    .CDOREADY_X0_Y1_D0               (o_if[1].ready),

    .CDIDATA_X0_Y2_D0                (i_if[2].data),
    .CDIVALID_X0_Y2_D0               (i_if[2].valid),
    .CDIREADY_X0_Y2_D0               (i_if[2].ready),
    .CDODATA_X0_Y2_D0                (o_if[2].data),
    .CDOVALID_X0_Y2_D0               (o_if[2].valid),
    .CDOREADY_X0_Y2_D0               (o_if[2].ready),

    .CDIDATA_X0_Y3_D0                (i_if[3].data),
    .CDIVALID_X0_Y3_D0               (i_if[3].valid),
    .CDIREADY_X0_Y3_D0               (i_if[3].ready),
    .CDODATA_X0_Y3_D0                (o_if[3].data),
    .CDOVALID_X0_Y3_D0               (o_if[3].valid),
    .CDOREADY_X0_Y3_D0               (o_if[3].ready),

    .CDIDATA_X0_Y4_D0                (i_if[4].data),
    .CDIVALID_X0_Y4_D0               (i_if[4].valid),
    .CDIREADY_X0_Y4_D0               (i_if[4].ready),
    .CDODATA_X0_Y4_D0                (o_if[4].data),
    .CDOVALID_X0_Y4_D0               (o_if[4].valid),
    .CDOREADY_X0_Y4_D0               (o_if[4].ready),

    .CDIDATA_X1_Y0_D0                (i_if[5].data),
    .CDIVALID_X1_Y0_D0               (i_if[5].valid),
    .CDIREADY_X1_Y0_D0               (i_if[5].ready),
    .CDODATA_X1_Y0_D0                (o_if[5].data),
    .CDOVALID_X1_Y0_D0               (o_if[5].valid),
    .CDOREADY_X1_Y0_D0               (o_if[5].ready),

    .CDIDATA_X1_Y1_D0                (i_if[6].data),
    .CDIVALID_X1_Y1_D0               (i_if[6].valid),
    .CDIREADY_X1_Y1_D0               (i_if[6].ready),
    .CDODATA_X1_Y1_D0                (o_if[6].data),
    .CDOVALID_X1_Y1_D0               (o_if[6].valid),
    .CDOREADY_X1_Y1_D0               (o_if[6].ready),

    .CDIDATA_X1_Y2_D0                (i_if[7].data),
    .CDIVALID_X1_Y2_D0               (i_if[7].valid),
    .CDIREADY_X1_Y2_D0               (i_if[7].ready),
    .CDODATA_X1_Y2_D0                (o_if[7].data),
    .CDOVALID_X1_Y2_D0               (o_if[7].valid),
    .CDOREADY_X1_Y2_D0               (o_if[7].ready),

    .CDIDATA_X1_Y3_D0                (i_if[8].data),
    .CDIVALID_X1_Y3_D0               (i_if[8].valid),
    .CDIREADY_X1_Y3_D0               (i_if[8].ready),
    .CDODATA_X1_Y3_D0                (o_if[8].data),
    .CDOVALID_X1_Y3_D0               (o_if[8].valid),
    .CDOREADY_X1_Y3_D0               (o_if[8].ready),

    .CDIDATA_X1_Y4_D0                (i_if[9].data),
    .CDIVALID_X1_Y4_D0               (i_if[9].valid),
    .CDIREADY_X1_Y4_D0               (i_if[9].ready),
    .CDODATA_X1_Y4_D0                (o_if[9].data),
    .CDOVALID_X1_Y4_D0               (o_if[9].valid),
    .CDOREADY_X1_Y4_D0               (o_if[9].ready),

    .CDIDATA_X2_Y1_D0                (i_if[11].data),
    .CDIVALID_X2_Y1_D0               (i_if[11].valid),
    .CDIREADY_X2_Y1_D0               (i_if[11].ready),
    .CDODATA_X2_Y1_D0                (o_if[11].data),
    .CDOVALID_X2_Y1_D0               (o_if[11].valid),
    .CDOREADY_X2_Y1_D0               (o_if[11].ready),

    .CDIDATA_X2_Y2_D0                (i_if[12].data),
    .CDIVALID_X2_Y2_D0               (i_if[12].valid),
    .CDIREADY_X2_Y2_D0               (i_if[12].ready),
    .CDODATA_X2_Y2_D0                (o_if[12].data),
    .CDOVALID_X2_Y2_D0               (o_if[12].valid),
    .CDOREADY_X2_Y2_D0               (o_if[12].ready),

    .CDIDATA_X2_Y3_D0                (i_if[13].data),
    .CDIVALID_X2_Y3_D0               (i_if[13].valid),
    .CDIREADY_X2_Y3_D0               (i_if[13].ready),
    .CDODATA_X2_Y3_D0                (o_if[13].data),
    .CDOVALID_X2_Y3_D0               (o_if[13].valid),
    .CDOREADY_X2_Y3_D0               (o_if[13].ready),

    .CDIDATA_X3_Y0_D0                (i_if[15].data),
    .CDIVALID_X3_Y0_D0               (i_if[15].valid),
    .CDIREADY_X3_Y0_D0               (i_if[15].ready),
    .CDODATA_X3_Y0_D0                (o_if[15].data),
    .CDOVALID_X3_Y0_D0               (o_if[15].valid),
    .CDOREADY_X3_Y0_D0               (o_if[15].ready),

    .CDIDATA_X3_Y1_D0                (i_if[16].data),
    .CDIVALID_X3_Y1_D0               (i_if[16].valid),
    .CDIREADY_X3_Y1_D0               (i_if[16].ready),
    .CDODATA_X3_Y1_D0                (o_if[16].data),
    .CDOVALID_X3_Y1_D0               (o_if[16].valid),
    .CDOREADY_X3_Y1_D0               (o_if[16].ready),

    .CDIDATA_X3_Y2_D0                (i_if[17].data),
    .CDIVALID_X3_Y2_D0               (i_if[17].valid),
    .CDIREADY_X3_Y2_D0               (i_if[17].ready),
    .CDODATA_X3_Y2_D0                (o_if[17].data),
    .CDOVALID_X3_Y2_D0               (o_if[17].valid),
    .CDOREADY_X3_Y2_D0               (o_if[17].ready),

    .CDIDATA_X3_Y3_D0                (i_if[18].data),
    .CDIVALID_X3_Y3_D0               (i_if[18].valid),
    .CDIREADY_X3_Y3_D0               (i_if[18].ready),
    .CDODATA_X3_Y3_D0                (o_if[18].data),
    .CDOVALID_X3_Y3_D0               (o_if[18].valid),
    .CDOREADY_X3_Y3_D0               (o_if[18].ready),

    .CDIDATA_X3_Y4_D0                (i_if[19].data),
    .CDIVALID_X3_Y4_D0               (i_if[19].valid),
    .CDIREADY_X3_Y4_D0               (i_if[19].ready),
    .CDODATA_X3_Y4_D0                (o_if[19].data),
    .CDOVALID_X3_Y4_D0               (o_if[19].valid),
    .CDOREADY_X3_Y4_D0               (o_if[19].ready),

    .CDIDATA_X4_Y0_D0                (i_if[20].data),
    .CDIVALID_X4_Y0_D0               (i_if[20].valid),
    .CDIREADY_X4_Y0_D0               (i_if[20].ready),
    .CDODATA_X4_Y0_D0                (o_if[20].data),
    .CDOVALID_X4_Y0_D0               (o_if[20].valid),
    .CDOREADY_X4_Y0_D0               (o_if[20].ready),

    .CDIDATA_X4_Y1_D0                (i_if[21].data),
    .CDIVALID_X4_Y1_D0               (i_if[21].valid),
    .CDIREADY_X4_Y1_D0               (i_if[21].ready),
    .CDODATA_X4_Y1_D0                (o_if[21].data),
    .CDOVALID_X4_Y1_D0               (o_if[21].valid),
    .CDOREADY_X4_Y1_D0               (o_if[21].ready),

    .CDIDATA_X4_Y2_D0                (i_if[22].data),
    .CDIVALID_X4_Y2_D0               (i_if[22].valid),
    .CDIREADY_X4_Y2_D0               (i_if[22].ready),
    .CDODATA_X4_Y2_D0                (o_if[22].data),
    .CDOVALID_X4_Y2_D0               (o_if[22].valid),
    .CDOREADY_X4_Y2_D0               (o_if[22].ready),

    .CDIDATA_X4_Y3_D0                (i_if[23].data),
    .CDIVALID_X4_Y3_D0               (i_if[23].valid),
    .CDIREADY_X4_Y3_D0               (i_if[23].ready),
    .CDODATA_X4_Y3_D0                (o_if[23].data),
    .CDOVALID_X4_Y3_D0               (o_if[23].valid),
    .CDOREADY_X4_Y3_D0               (o_if[23].ready),

    .CDIDATA_X4_Y4_D0                (i_if[24].data),
    .CDIVALID_X4_Y4_D0               (i_if[24].valid),
    .CDIREADY_X4_Y4_D0               (i_if[24].ready),
    .CDODATA_X4_Y4_D0                (o_if[24].data),
    .CDOVALID_X4_Y4_D0               (o_if[24].valid),
    .CDOREADY_X4_Y4_D0               (o_if[24].ready),

    .CDIDATA_X0_Y0_D1                (i_if[25].data),
    .CDIVALID_X0_Y0_D1               (i_if[25].valid),
    .CDIREADY_X0_Y0_D1               (i_if[25].ready),
    .CDODATA_X0_Y0_D1                (o_if[25].data),
    .CDOVALID_X0_Y0_D1               (o_if[25].valid),
    .CDOREADY_X0_Y0_D1               (o_if[25].ready),

    .CDIDATA_X0_Y1_D1                (i_if[26].data),
    .CDIVALID_X0_Y1_D1               (i_if[26].valid),
    .CDIREADY_X0_Y1_D1               (i_if[26].ready),
    .CDODATA_X0_Y1_D1                (o_if[26].data),
    .CDOVALID_X0_Y1_D1               (o_if[26].valid),
    .CDOREADY_X0_Y1_D1               (o_if[26].ready),

    .CDIDATA_X0_Y2_D1                (i_if[27].data),
    .CDIVALID_X0_Y2_D1               (i_if[27].valid),
    .CDIREADY_X0_Y2_D1               (i_if[27].ready),
    .CDODATA_X0_Y2_D1                (o_if[27].data),
    .CDOVALID_X0_Y2_D1               (o_if[27].valid),
    .CDOREADY_X0_Y2_D1               (o_if[27].ready),

    .CDIDATA_X0_Y3_D1                (i_if[28].data),
    .CDIVALID_X0_Y3_D1               (i_if[28].valid),
    .CDIREADY_X0_Y3_D1               (i_if[28].ready),
    .CDODATA_X0_Y3_D1                (o_if[28].data),
    .CDOVALID_X0_Y3_D1               (o_if[28].valid),
    .CDOREADY_X0_Y3_D1               (o_if[28].ready),

    .CDIDATA_X0_Y4_D1                (i_if[29].data),
    .CDIVALID_X0_Y4_D1               (i_if[29].valid),
    .CDIREADY_X0_Y4_D1               (i_if[29].ready),
    .CDODATA_X0_Y4_D1                (o_if[29].data),
    .CDOVALID_X0_Y4_D1               (o_if[29].valid),
    .CDOREADY_X0_Y4_D1               (o_if[29].ready),

    .CDIDATA_X1_Y0_D1                (i_if[30].data),
    .CDIVALID_X1_Y0_D1               (i_if[30].valid),
    .CDIREADY_X1_Y0_D1               (i_if[30].ready),
    .CDODATA_X1_Y0_D1                (o_if[30].data),
    .CDOVALID_X1_Y0_D1               (o_if[30].valid),
    .CDOREADY_X1_Y0_D1               (o_if[30].ready),

    .CDIDATA_X1_Y1_D1                (i_if[31].data),
    .CDIVALID_X1_Y1_D1               (i_if[31].valid),
    .CDIREADY_X1_Y1_D1               (i_if[31].ready),
    .CDODATA_X1_Y1_D1                (o_if[31].data),
    .CDOVALID_X1_Y1_D1               (o_if[31].valid),
    .CDOREADY_X1_Y1_D1               (o_if[31].ready),

    .CDIDATA_X1_Y2_D1                (i_if[32].data),
    .CDIVALID_X1_Y2_D1               (i_if[32].valid),
    .CDIREADY_X1_Y2_D1               (i_if[32].ready),
    .CDODATA_X1_Y2_D1                (o_if[32].data),
    .CDOVALID_X1_Y2_D1               (o_if[32].valid),
    .CDOREADY_X1_Y2_D1               (o_if[32].ready),

    .CDIDATA_X1_Y3_D1                (i_if[33].data),
    .CDIVALID_X1_Y3_D1               (i_if[33].valid),
    .CDIREADY_X1_Y3_D1               (i_if[33].ready),
    .CDODATA_X1_Y3_D1                (o_if[33].data),
    .CDOVALID_X1_Y3_D1               (o_if[33].valid),
    .CDOREADY_X1_Y3_D1               (o_if[33].ready),

    .CDIDATA_X1_Y4_D1                (i_if[34].data),
    .CDIVALID_X1_Y4_D1               (i_if[34].valid),
    .CDIREADY_X1_Y4_D1               (i_if[34].ready),
    .CDODATA_X1_Y4_D1                (o_if[34].data),
    .CDOVALID_X1_Y4_D1               (o_if[34].valid),
    .CDOREADY_X1_Y4_D1               (o_if[34].ready),

    .CDIDATA_X2_Y1_D1                (i_if[36].data),
    .CDIVALID_X2_Y1_D1               (i_if[36].valid),
    .CDIREADY_X2_Y1_D1               (i_if[36].ready),
    .CDODATA_X2_Y1_D1                (o_if[36].data),
    .CDOVALID_X2_Y1_D1               (o_if[36].valid),
    .CDOREADY_X2_Y1_D1               (o_if[36].ready),

    .CDIDATA_X2_Y2_D1                (i_if[37].data),
    .CDIVALID_X2_Y2_D1               (i_if[37].valid),
    .CDIREADY_X2_Y2_D1               (i_if[37].ready),
    .CDODATA_X2_Y2_D1                (o_if[37].data),
    .CDOVALID_X2_Y2_D1               (o_if[37].valid),
    .CDOREADY_X2_Y2_D1               (o_if[37].ready),

    .CDIDATA_X2_Y3_D1                (i_if[38].data),
    .CDIVALID_X2_Y3_D1               (i_if[38].valid),
    .CDIREADY_X2_Y3_D1               (i_if[38].ready),
    .CDODATA_X2_Y3_D1                (o_if[38].data),
    .CDOVALID_X2_Y3_D1               (o_if[38].valid),
    .CDOREADY_X2_Y3_D1               (o_if[38].ready),

    .CDIDATA_X3_Y0_D1                (i_if[40].data),
    .CDIVALID_X3_Y0_D1               (i_if[40].valid),
    .CDIREADY_X3_Y0_D1               (i_if[40].ready),
    .CDODATA_X3_Y0_D1                (o_if[40].data),
    .CDOVALID_X3_Y0_D1               (o_if[40].valid),
    .CDOREADY_X3_Y0_D1               (o_if[40].ready),

    .CDIDATA_X3_Y1_D1                (i_if[41].data),
    .CDIVALID_X3_Y1_D1               (i_if[41].valid),
    .CDIREADY_X3_Y1_D1               (i_if[41].ready),
    .CDODATA_X3_Y1_D1                (o_if[41].data),
    .CDOVALID_X3_Y1_D1               (o_if[41].valid),
    .CDOREADY_X3_Y1_D1               (o_if[41].ready),

    .CDIDATA_X3_Y2_D1                (i_if[42].data),
    .CDIVALID_X3_Y2_D1               (i_if[42].valid),
    .CDIREADY_X3_Y2_D1               (i_if[42].ready),
    .CDODATA_X3_Y2_D1                (o_if[42].data),
    .CDOVALID_X3_Y2_D1               (o_if[42].valid),
    .CDOREADY_X3_Y2_D1               (o_if[42].ready),

    .CDIDATA_X3_Y3_D1                (i_if[43].data),
    .CDIVALID_X3_Y3_D1               (i_if[43].valid),
    .CDIREADY_X3_Y3_D1               (i_if[43].ready),
    .CDODATA_X3_Y3_D1                (o_if[43].data),
    .CDOVALID_X3_Y3_D1               (o_if[43].valid),
    .CDOREADY_X3_Y3_D1               (o_if[43].ready),

    .CDIDATA_X3_Y4_D1                (i_if[44].data),
    .CDIVALID_X3_Y4_D1               (i_if[44].valid),
    .CDIREADY_X3_Y4_D1               (i_if[44].ready),
    .CDODATA_X3_Y4_D1                (o_if[44].data),
    .CDOVALID_X3_Y4_D1               (o_if[44].valid),
    .CDOREADY_X3_Y4_D1               (o_if[44].ready),

    .CDIDATA_X4_Y0_D1                (i_if[45].data),
    .CDIVALID_X4_Y0_D1               (i_if[45].valid),
    .CDIREADY_X4_Y0_D1               (i_if[45].ready),
    .CDODATA_X4_Y0_D1                (o_if[45].data),
    .CDOVALID_X4_Y0_D1               (o_if[45].valid),
    .CDOREADY_X4_Y0_D1               (o_if[45].ready),

    .CDIDATA_X4_Y1_D1                (i_if[46].data),
    .CDIVALID_X4_Y1_D1               (i_if[46].valid),
    .CDIREADY_X4_Y1_D1               (i_if[46].ready),
    .CDODATA_X4_Y1_D1                (o_if[46].data),
    .CDOVALID_X4_Y1_D1               (o_if[46].valid),
    .CDOREADY_X4_Y1_D1               (o_if[46].ready),

    .CDIDATA_X4_Y2_D1                (i_if[47].data),
    .CDIVALID_X4_Y2_D1               (i_if[47].valid),
    .CDIREADY_X4_Y2_D1               (i_if[47].ready),
    .CDODATA_X4_Y2_D1                (o_if[47].data),
    .CDOVALID_X4_Y2_D1               (o_if[47].valid),
    .CDOREADY_X4_Y2_D1               (o_if[47].ready),

    .CDIDATA_X4_Y3_D1                (i_if[48].data),
    .CDIVALID_X4_Y3_D1               (i_if[48].valid),
    .CDIREADY_X4_Y3_D1               (i_if[48].ready),
    .CDODATA_X4_Y3_D1                (o_if[48].data),
    .CDOVALID_X4_Y3_D1               (o_if[48].valid),
    .CDOREADY_X4_Y3_D1               (o_if[48].ready),

    .CDIDATA_X4_Y4_D1                (i_if[49].data),
    .CDIVALID_X4_Y4_D1               (i_if[49].valid),
    .CDIREADY_X4_Y4_D1               (i_if[49].ready),
    .CDODATA_X4_Y4_D1                (o_if[49].data),
    .CDOVALID_X4_Y4_D1               (o_if[49].valid),
    .CDOREADY_X4_Y4_D1               (o_if[49].ready),

    .CDIDATA_X0_Y0_D2                (i_if[50].data),
    .CDIVALID_X0_Y0_D2               (i_if[50].valid),
    .CDIREADY_X0_Y0_D2               (i_if[50].ready),
    .CDODATA_X0_Y0_D2                (o_if[50].data),
    .CDOVALID_X0_Y0_D2               (o_if[50].valid),
    .CDOREADY_X0_Y0_D2               (o_if[50].ready),

    .CDIDATA_X0_Y1_D2                (i_if[51].data),
    .CDIVALID_X0_Y1_D2               (i_if[51].valid),
    .CDIREADY_X0_Y1_D2               (i_if[51].ready),
    .CDODATA_X0_Y1_D2                (o_if[51].data),
    .CDOVALID_X0_Y1_D2               (o_if[51].valid),
    .CDOREADY_X0_Y1_D2               (o_if[51].ready),

    .CDIDATA_X0_Y2_D2                (i_if[52].data),
    .CDIVALID_X0_Y2_D2               (i_if[52].valid),
    .CDIREADY_X0_Y2_D2               (i_if[52].ready),
    .CDODATA_X0_Y2_D2                (o_if[52].data),
    .CDOVALID_X0_Y2_D2               (o_if[52].valid),
    .CDOREADY_X0_Y2_D2               (o_if[52].ready),

    .CDIDATA_X0_Y3_D2                (i_if[53].data),
    .CDIVALID_X0_Y3_D2               (i_if[53].valid),
    .CDIREADY_X0_Y3_D2               (i_if[53].ready),
    .CDODATA_X0_Y3_D2                (o_if[53].data),
    .CDOVALID_X0_Y3_D2               (o_if[53].valid),
    .CDOREADY_X0_Y3_D2               (o_if[53].ready),

    .CDIDATA_X0_Y4_D2                (i_if[54].data),
    .CDIVALID_X0_Y4_D2               (i_if[54].valid),
    .CDIREADY_X0_Y4_D2               (i_if[54].ready),
    .CDODATA_X0_Y4_D2                (o_if[54].data),
    .CDOVALID_X0_Y4_D2               (o_if[54].valid),
    .CDOREADY_X0_Y4_D2               (o_if[54].ready),

    .CDIDATA_X1_Y0_D2                (i_if[55].data),
    .CDIVALID_X1_Y0_D2               (i_if[55].valid),
    .CDIREADY_X1_Y0_D2               (i_if[55].ready),
    .CDODATA_X1_Y0_D2                (o_if[55].data),
    .CDOVALID_X1_Y0_D2               (o_if[55].valid),
    .CDOREADY_X1_Y0_D2               (o_if[55].ready),

    .CDIDATA_X1_Y1_D2                (i_if[56].data),
    .CDIVALID_X1_Y1_D2               (i_if[56].valid),
    .CDIREADY_X1_Y1_D2               (i_if[56].ready),
    .CDODATA_X1_Y1_D2                (o_if[56].data),
    .CDOVALID_X1_Y1_D2               (o_if[56].valid),
    .CDOREADY_X1_Y1_D2               (o_if[56].ready),

    .CDIDATA_X1_Y2_D2                (i_if[57].data),
    .CDIVALID_X1_Y2_D2               (i_if[57].valid),
    .CDIREADY_X1_Y2_D2               (i_if[57].ready),
    .CDODATA_X1_Y2_D2                (o_if[57].data),
    .CDOVALID_X1_Y2_D2               (o_if[57].valid),
    .CDOREADY_X1_Y2_D2               (o_if[57].ready),

    .CDIDATA_X1_Y3_D2                (i_if[58].data),
    .CDIVALID_X1_Y3_D2               (i_if[58].valid),
    .CDIREADY_X1_Y3_D2               (i_if[58].ready),
    .CDODATA_X1_Y3_D2                (o_if[58].data),
    .CDOVALID_X1_Y3_D2               (o_if[58].valid),
    .CDOREADY_X1_Y3_D2               (o_if[58].ready),

    .CDIDATA_X1_Y4_D2                (i_if[59].data),
    .CDIVALID_X1_Y4_D2               (i_if[59].valid),
    .CDIREADY_X1_Y4_D2               (i_if[59].ready),
    .CDODATA_X1_Y4_D2                (o_if[59].data),
    .CDOVALID_X1_Y4_D2               (o_if[59].valid),
    .CDOREADY_X1_Y4_D2               (o_if[59].ready),

    .CDIDATA_X2_Y1_D2                (i_if[61].data),
    .CDIVALID_X2_Y1_D2               (i_if[61].valid),
    .CDIREADY_X2_Y1_D2               (i_if[61].ready),
    .CDODATA_X2_Y1_D2                (o_if[61].data),
    .CDOVALID_X2_Y1_D2               (o_if[61].valid),
    .CDOREADY_X2_Y1_D2               (o_if[61].ready),

    .CDIDATA_X2_Y2_D2                (i_if[62].data),
    .CDIVALID_X2_Y2_D2               (i_if[62].valid),
    .CDIREADY_X2_Y2_D2               (i_if[62].ready),
    .CDODATA_X2_Y2_D2                (o_if[62].data),
    .CDOVALID_X2_Y2_D2               (o_if[62].valid),
    .CDOREADY_X2_Y2_D2               (o_if[62].ready),

    .CDIDATA_X2_Y3_D2                (i_if[63].data),
    .CDIVALID_X2_Y3_D2               (i_if[63].valid),
    .CDIREADY_X2_Y3_D2               (i_if[63].ready),
    .CDODATA_X2_Y3_D2                (o_if[63].data),
    .CDOVALID_X2_Y3_D2               (o_if[63].valid),
    .CDOREADY_X2_Y3_D2               (o_if[63].ready),

    .CDIDATA_X3_Y0_D2                (i_if[65].data),
    .CDIVALID_X3_Y0_D2               (i_if[65].valid),
    .CDIREADY_X3_Y0_D2               (i_if[65].ready),
    .CDODATA_X3_Y0_D2                (o_if[65].data),
    .CDOVALID_X3_Y0_D2               (o_if[65].valid),
    .CDOREADY_X3_Y0_D2               (o_if[65].ready),

    .CDIDATA_X3_Y1_D2                (i_if[66].data),
    .CDIVALID_X3_Y1_D2               (i_if[66].valid),
    .CDIREADY_X3_Y1_D2               (i_if[66].ready),
    .CDODATA_X3_Y1_D2                (o_if[66].data),
    .CDOVALID_X3_Y1_D2               (o_if[66].valid),
    .CDOREADY_X3_Y1_D2               (o_if[66].ready),

    .CDIDATA_X3_Y2_D2                (i_if[67].data),
    .CDIVALID_X3_Y2_D2               (i_if[67].valid),
    .CDIREADY_X3_Y2_D2               (i_if[67].ready),
    .CDODATA_X3_Y2_D2                (o_if[67].data),
    .CDOVALID_X3_Y2_D2               (o_if[67].valid),
    .CDOREADY_X3_Y2_D2               (o_if[67].ready),

    .CDIDATA_X3_Y3_D2                (i_if[68].data),
    .CDIVALID_X3_Y3_D2               (i_if[68].valid),
    .CDIREADY_X3_Y3_D2               (i_if[68].ready),
    .CDODATA_X3_Y3_D2                (o_if[68].data),
    .CDOVALID_X3_Y3_D2               (o_if[68].valid),
    .CDOREADY_X3_Y3_D2               (o_if[68].ready),

    .CDIDATA_X3_Y4_D2                (i_if[69].data),
    .CDIVALID_X3_Y4_D2               (i_if[69].valid),
    .CDIREADY_X3_Y4_D2               (i_if[69].ready),
    .CDODATA_X3_Y4_D2                (o_if[69].data),
    .CDOVALID_X3_Y4_D2               (o_if[69].valid),
    .CDOREADY_X3_Y4_D2               (o_if[69].ready),

    .CDIDATA_X4_Y0_D2                (i_if[70].data),
    .CDIVALID_X4_Y0_D2               (i_if[70].valid),
    .CDIREADY_X4_Y0_D2               (i_if[70].ready),
    .CDODATA_X4_Y0_D2                (o_if[70].data),
    .CDOVALID_X4_Y0_D2               (o_if[70].valid),
    .CDOREADY_X4_Y0_D2               (o_if[70].ready),

    .CDIDATA_X4_Y1_D2                (i_if[71].data),
    .CDIVALID_X4_Y1_D2               (i_if[71].valid),
    .CDIREADY_X4_Y1_D2               (i_if[71].ready),
    .CDODATA_X4_Y1_D2                (o_if[71].data),
    .CDOVALID_X4_Y1_D2               (o_if[71].valid),
    .CDOREADY_X4_Y1_D2               (o_if[71].ready),

    .CDIDATA_X4_Y2_D2                (i_if[72].data),
    .CDIVALID_X4_Y2_D2               (i_if[72].valid),
    .CDIREADY_X4_Y2_D2               (i_if[72].ready),
    .CDODATA_X4_Y2_D2                (o_if[72].data),
    .CDOVALID_X4_Y2_D2               (o_if[72].valid),
    .CDOREADY_X4_Y2_D2               (o_if[72].ready),

    .CDIDATA_X4_Y3_D2                (i_if[73].data),
    .CDIVALID_X4_Y3_D2               (i_if[73].valid),
    .CDIREADY_X4_Y3_D2               (i_if[73].ready),
    .CDODATA_X4_Y3_D2                (o_if[73].data),
    .CDOVALID_X4_Y3_D2               (o_if[73].valid),
    .CDOREADY_X4_Y3_D2               (o_if[73].ready),

    .CDIDATA_X4_Y4_D2                (i_if[74].data),
    .CDIVALID_X4_Y4_D2               (i_if[74].valid),
    .CDIREADY_X4_Y4_D2               (i_if[74].ready),
    .CDODATA_X4_Y4_D2                (o_if[74].data),
    .CDOVALID_X4_Y4_D2               (o_if[74].valid),
    .CDOREADY_X4_Y4_D2               (o_if[74].ready)
);

initial
begin
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[0].drv","vif",i_if[0]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[0].mon","vif",o_if[0]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[1].drv","vif",i_if[1]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[1].mon","vif",o_if[1]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[2].drv","vif",i_if[2]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[2].mon","vif",o_if[2]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[3].drv","vif",i_if[3]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[3].mon","vif",o_if[3]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[4].drv","vif",i_if[4]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[4].mon","vif",o_if[4]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[5].drv","vif",i_if[5]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[5].mon","vif",o_if[5]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[6].drv","vif",i_if[6]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[6].mon","vif",o_if[6]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[7].drv","vif",i_if[7]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[7].mon","vif",o_if[7]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[8].drv","vif",i_if[8]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[8].mon","vif",o_if[8]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[9].drv","vif",i_if[9]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[9].mon","vif",o_if[9]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[11].drv","vif",i_if[11]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[11].mon","vif",o_if[11]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[12].drv","vif",i_if[12]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[12].mon","vif",o_if[12]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[13].drv","vif",i_if[13]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[13].mon","vif",o_if[13]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[15].drv","vif",i_if[15]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[15].mon","vif",o_if[15]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[16].drv","vif",i_if[16]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[16].mon","vif",o_if[16]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[17].drv","vif",i_if[17]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[17].mon","vif",o_if[17]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[18].drv","vif",i_if[18]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[18].mon","vif",o_if[18]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[19].drv","vif",i_if[19]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[19].mon","vif",o_if[19]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[20].drv","vif",i_if[20]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[20].mon","vif",o_if[20]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[21].drv","vif",i_if[21]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[21].mon","vif",o_if[21]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[22].drv","vif",i_if[22]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[22].mon","vif",o_if[22]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[23].drv","vif",i_if[23]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[23].mon","vif",o_if[23]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[24].drv","vif",i_if[24]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[24].mon","vif",o_if[24]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[25].drv","vif",i_if[25]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[25].mon","vif",o_if[25]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[26].drv","vif",i_if[26]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[26].mon","vif",o_if[26]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[27].drv","vif",i_if[27]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[27].mon","vif",o_if[27]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[28].drv","vif",i_if[28]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[28].mon","vif",o_if[28]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[29].drv","vif",i_if[29]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[29].mon","vif",o_if[29]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[30].drv","vif",i_if[30]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[30].mon","vif",o_if[30]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[31].drv","vif",i_if[31]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[31].mon","vif",o_if[31]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[32].drv","vif",i_if[32]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[32].mon","vif",o_if[32]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[33].drv","vif",i_if[33]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[33].mon","vif",o_if[33]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[34].drv","vif",i_if[34]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[34].mon","vif",o_if[34]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[36].drv","vif",i_if[36]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[36].mon","vif",o_if[36]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[37].drv","vif",i_if[37]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[37].mon","vif",o_if[37]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[38].drv","vif",i_if[38]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[38].mon","vif",o_if[38]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[40].drv","vif",i_if[40]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[40].mon","vif",o_if[40]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[41].drv","vif",i_if[41]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[41].mon","vif",o_if[41]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[42].drv","vif",i_if[42]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[42].mon","vif",o_if[42]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[43].drv","vif",i_if[43]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[43].mon","vif",o_if[43]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[44].drv","vif",i_if[44]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[44].mon","vif",o_if[44]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[45].drv","vif",i_if[45]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[45].mon","vif",o_if[45]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[46].drv","vif",i_if[46]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[46].mon","vif",o_if[46]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[47].drv","vif",i_if[47]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[47].mon","vif",o_if[47]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[48].drv","vif",i_if[48]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[48].mon","vif",o_if[48]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[49].drv","vif",i_if[49]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[49].mon","vif",o_if[49]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[50].drv","vif",i_if[50]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[50].mon","vif",o_if[50]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[51].drv","vif",i_if[51]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[51].mon","vif",o_if[51]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[52].drv","vif",i_if[52]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[52].mon","vif",o_if[52]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[53].drv","vif",i_if[53]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[53].mon","vif",o_if[53]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[54].drv","vif",i_if[54]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[54].mon","vif",o_if[54]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[55].drv","vif",i_if[55]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[55].mon","vif",o_if[55]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[56].drv","vif",i_if[56]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[56].mon","vif",o_if[56]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[57].drv","vif",i_if[57]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[57].mon","vif",o_if[57]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[58].drv","vif",i_if[58]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[58].mon","vif",o_if[58]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[59].drv","vif",i_if[59]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[59].mon","vif",o_if[59]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[61].drv","vif",i_if[61]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[61].mon","vif",o_if[61]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[62].drv","vif",i_if[62]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[62].mon","vif",o_if[62]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[63].drv","vif",i_if[63]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[63].mon","vif",o_if[63]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[65].drv","vif",i_if[65]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[65].mon","vif",o_if[65]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[66].drv","vif",i_if[66]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[66].mon","vif",o_if[66]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[67].drv","vif",i_if[67]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[67].mon","vif",o_if[67]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[68].drv","vif",i_if[68]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[68].mon","vif",o_if[68]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[69].drv","vif",i_if[69]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[69].mon","vif",o_if[69]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[70].drv","vif",i_if[70]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[70].mon","vif",o_if[70]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[71].drv","vif",i_if[71]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[71].mon","vif",o_if[71]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[72].drv","vif",i_if[72]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[72].mon","vif",o_if[72]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[73].drv","vif",i_if[73]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[73].mon","vif",o_if[73]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.i_agt[74].drv","vif",i_if[74]);
    uvm_config_db #(virtual cibd_if)::set(null,"uvm_test_top.env.o_agt[74].mon","vif",o_if[74]);
end

initial
begin
    run_test("nop_case0");
end

initial
begin
    clk_d = 0;
    forever
    begin
        #(`CD_CYCLE/2) clk_d = ~clk_d;
    end
end

initial
begin
    clk_p = 0;
    forever
    begin
        #(`CP_CYCLE/2) clk_p = ~clk_p;
    end
end

initial
begin
    rstn = 1'b0;
    #73;
    rstn = 1'b1;
end

endmodule