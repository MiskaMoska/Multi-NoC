interface cibd_if(input clk,input rstn);

    logic [129:0] data;
    logic valid,ready;
    
endinterface