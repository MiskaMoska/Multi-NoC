//Network on Chip
//Width: 5
//Height:5
`include "param.vh"

module NoD #(
    parameter NODID = 0
)(
    input       wire                                CDCLK,
    input       wire                                CDRESETn,
    
    //router0
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X0_Y0,
    input       wire                                CDIVALID_X0_Y0,
    output      wire                                CDIREADY_X0_Y0,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X0_Y0,
    output      wire                                CDOVALID_X0_Y0,
    input       wire                                CDOREADY_X0_Y0,

    //router1
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X0_Y1,
    input       wire                                CDIVALID_X0_Y1,
    output      wire                                CDIREADY_X0_Y1,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X0_Y1,
    output      wire                                CDOVALID_X0_Y1,
    input       wire                                CDOREADY_X0_Y1,

    //router2
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X0_Y2,
    input       wire                                CDIVALID_X0_Y2,
    output      wire                                CDIREADY_X0_Y2,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X0_Y2,
    output      wire                                CDOVALID_X0_Y2,
    input       wire                                CDOREADY_X0_Y2,

    //router3
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X0_Y3,
    input       wire                                CDIVALID_X0_Y3,
    output      wire                                CDIREADY_X0_Y3,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X0_Y3,
    output      wire                                CDOVALID_X0_Y3,
    input       wire                                CDOREADY_X0_Y3,

    //router4
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X0_Y4,
    input       wire                                CDIVALID_X0_Y4,
    output      wire                                CDIREADY_X0_Y4,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X0_Y4,
    output      wire                                CDOVALID_X0_Y4,
    input       wire                                CDOREADY_X0_Y4,

    //router5
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X1_Y0,
    input       wire                                CDIVALID_X1_Y0,
    output      wire                                CDIREADY_X1_Y0,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X1_Y0,
    output      wire                                CDOVALID_X1_Y0,
    input       wire                                CDOREADY_X1_Y0,

    //router6
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X1_Y1,
    input       wire                                CDIVALID_X1_Y1,
    output      wire                                CDIREADY_X1_Y1,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X1_Y1,
    output      wire                                CDOVALID_X1_Y1,
    input       wire                                CDOREADY_X1_Y1,

    //router7
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X1_Y2,
    input       wire                                CDIVALID_X1_Y2,
    output      wire                                CDIREADY_X1_Y2,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X1_Y2,
    output      wire                                CDOVALID_X1_Y2,
    input       wire                                CDOREADY_X1_Y2,

    //router8
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X1_Y3,
    input       wire                                CDIVALID_X1_Y3,
    output      wire                                CDIREADY_X1_Y3,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X1_Y3,
    output      wire                                CDOVALID_X1_Y3,
    input       wire                                CDOREADY_X1_Y3,

    //router9
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X1_Y4,
    input       wire                                CDIVALID_X1_Y4,
    output      wire                                CDIREADY_X1_Y4,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X1_Y4,
    output      wire                                CDOVALID_X1_Y4,
    input       wire                                CDOREADY_X1_Y4,

    //router10
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X2_Y0,
    input       wire                                CDIVALID_X2_Y0,
    output      wire                                CDIREADY_X2_Y0,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X2_Y0,
    output      wire                                CDOVALID_X2_Y0,
    input       wire                                CDOREADY_X2_Y0,

    //router11
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X2_Y1,
    input       wire                                CDIVALID_X2_Y1,
    output      wire                                CDIREADY_X2_Y1,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X2_Y1,
    output      wire                                CDOVALID_X2_Y1,
    input       wire                                CDOREADY_X2_Y1,

    //router12
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X2_Y2,
    input       wire                                CDIVALID_X2_Y2,
    output      wire                                CDIREADY_X2_Y2,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X2_Y2,
    output      wire                                CDOVALID_X2_Y2,
    input       wire                                CDOREADY_X2_Y2,

    //router13
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X2_Y3,
    input       wire                                CDIVALID_X2_Y3,
    output      wire                                CDIREADY_X2_Y3,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X2_Y3,
    output      wire                                CDOVALID_X2_Y3,
    input       wire                                CDOREADY_X2_Y3,

    //router14
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X2_Y4,
    input       wire                                CDIVALID_X2_Y4,
    output      wire                                CDIREADY_X2_Y4,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X2_Y4,
    output      wire                                CDOVALID_X2_Y4,
    input       wire                                CDOREADY_X2_Y4,

    //router15
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X3_Y0,
    input       wire                                CDIVALID_X3_Y0,
    output      wire                                CDIREADY_X3_Y0,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X3_Y0,
    output      wire                                CDOVALID_X3_Y0,
    input       wire                                CDOREADY_X3_Y0,

    //router16
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X3_Y1,
    input       wire                                CDIVALID_X3_Y1,
    output      wire                                CDIREADY_X3_Y1,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X3_Y1,
    output      wire                                CDOVALID_X3_Y1,
    input       wire                                CDOREADY_X3_Y1,

    //router17
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X3_Y2,
    input       wire                                CDIVALID_X3_Y2,
    output      wire                                CDIREADY_X3_Y2,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X3_Y2,
    output      wire                                CDOVALID_X3_Y2,
    input       wire                                CDOREADY_X3_Y2,

    //router18
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X3_Y3,
    input       wire                                CDIVALID_X3_Y3,
    output      wire                                CDIREADY_X3_Y3,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X3_Y3,
    output      wire                                CDOVALID_X3_Y3,
    input       wire                                CDOREADY_X3_Y3,

    //router19
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X3_Y4,
    input       wire                                CDIVALID_X3_Y4,
    output      wire                                CDIREADY_X3_Y4,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X3_Y4,
    output      wire                                CDOVALID_X3_Y4,
    input       wire                                CDOREADY_X3_Y4,

    //router20
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X4_Y0,
    input       wire                                CDIVALID_X4_Y0,
    output      wire                                CDIREADY_X4_Y0,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X4_Y0,
    output      wire                                CDOVALID_X4_Y0,
    input       wire                                CDOREADY_X4_Y0,

    //router21
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X4_Y1,
    input       wire                                CDIVALID_X4_Y1,
    output      wire                                CDIREADY_X4_Y1,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X4_Y1,
    output      wire                                CDOVALID_X4_Y1,
    input       wire                                CDOREADY_X4_Y1,

    //router22
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X4_Y2,
    input       wire                                CDIVALID_X4_Y2,
    output      wire                                CDIREADY_X4_Y2,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X4_Y2,
    output      wire                                CDOVALID_X4_Y2,
    input       wire                                CDOREADY_X4_Y2,

    //router23
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X4_Y3,
    input       wire                                CDIVALID_X4_Y3,
    output      wire                                CDIREADY_X4_Y3,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X4_Y3,
    output      wire                                CDOVALID_X4_Y3,
    input       wire                                CDOREADY_X4_Y3,

    //router24
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X4_Y4,
    input       wire                                CDIVALID_X4_Y4,
    output      wire                                CDIREADY_X4_Y4,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X4_Y4,
    output      wire                                CDOVALID_X4_Y4,
    input       wire                                CDOREADY_X4_Y4
);

//horizontal signals
wire    [`DATA_WIDTH-1:0]   data_0_to_1,	data_1_to_0;
wire                        valid_0_to_1,	valid_1_to_0;
wire                        ready_0_to_1,	ready_1_to_0;
wire    [`DATA_WIDTH-1:0]   data_1_to_2,	data_2_to_1;
wire                        valid_1_to_2,	valid_2_to_1;
wire                        ready_1_to_2,	ready_2_to_1;
wire    [`DATA_WIDTH-1:0]   data_2_to_3,	data_3_to_2;
wire                        valid_2_to_3,	valid_3_to_2;
wire                        ready_2_to_3,	ready_3_to_2;
wire    [`DATA_WIDTH-1:0]   data_3_to_4,	data_4_to_3;
wire                        valid_3_to_4,	valid_4_to_3;
wire                        ready_3_to_4,	ready_4_to_3;
wire    [`DATA_WIDTH-1:0]   data_5_to_6,	data_6_to_5;
wire                        valid_5_to_6,	valid_6_to_5;
wire                        ready_5_to_6,	ready_6_to_5;
wire    [`DATA_WIDTH-1:0]   data_6_to_7,	data_7_to_6;
wire                        valid_6_to_7,	valid_7_to_6;
wire                        ready_6_to_7,	ready_7_to_6;
wire    [`DATA_WIDTH-1:0]   data_7_to_8,	data_8_to_7;
wire                        valid_7_to_8,	valid_8_to_7;
wire                        ready_7_to_8,	ready_8_to_7;
wire    [`DATA_WIDTH-1:0]   data_8_to_9,	data_9_to_8;
wire                        valid_8_to_9,	valid_9_to_8;
wire                        ready_8_to_9,	ready_9_to_8;
wire    [`DATA_WIDTH-1:0]   data_10_to_11,	data_11_to_10;
wire                        valid_10_to_11,	valid_11_to_10;
wire                        ready_10_to_11,	ready_11_to_10;
wire    [`DATA_WIDTH-1:0]   data_11_to_12,	data_12_to_11;
wire                        valid_11_to_12,	valid_12_to_11;
wire                        ready_11_to_12,	ready_12_to_11;
wire    [`DATA_WIDTH-1:0]   data_12_to_13,	data_13_to_12;
wire                        valid_12_to_13,	valid_13_to_12;
wire                        ready_12_to_13,	ready_13_to_12;
wire    [`DATA_WIDTH-1:0]   data_13_to_14,	data_14_to_13;
wire                        valid_13_to_14,	valid_14_to_13;
wire                        ready_13_to_14,	ready_14_to_13;
wire    [`DATA_WIDTH-1:0]   data_15_to_16,	data_16_to_15;
wire                        valid_15_to_16,	valid_16_to_15;
wire                        ready_15_to_16,	ready_16_to_15;
wire    [`DATA_WIDTH-1:0]   data_16_to_17,	data_17_to_16;
wire                        valid_16_to_17,	valid_17_to_16;
wire                        ready_16_to_17,	ready_17_to_16;
wire    [`DATA_WIDTH-1:0]   data_17_to_18,	data_18_to_17;
wire                        valid_17_to_18,	valid_18_to_17;
wire                        ready_17_to_18,	ready_18_to_17;
wire    [`DATA_WIDTH-1:0]   data_18_to_19,	data_19_to_18;
wire                        valid_18_to_19,	valid_19_to_18;
wire                        ready_18_to_19,	ready_19_to_18;
wire    [`DATA_WIDTH-1:0]   data_20_to_21,	data_21_to_20;
wire                        valid_20_to_21,	valid_21_to_20;
wire                        ready_20_to_21,	ready_21_to_20;
wire    [`DATA_WIDTH-1:0]   data_21_to_22,	data_22_to_21;
wire                        valid_21_to_22,	valid_22_to_21;
wire                        ready_21_to_22,	ready_22_to_21;
wire    [`DATA_WIDTH-1:0]   data_22_to_23,	data_23_to_22;
wire                        valid_22_to_23,	valid_23_to_22;
wire                        ready_22_to_23,	ready_23_to_22;
wire    [`DATA_WIDTH-1:0]   data_23_to_24,	data_24_to_23;
wire                        valid_23_to_24,	valid_24_to_23;
wire                        ready_23_to_24,	ready_24_to_23;

//vertical signals
wire    [`DATA_WIDTH-1:0]   data_0_to_5,	data_5_to_0;
wire                        valid_0_to_5,	valid_5_to_0;
wire                        ready_0_to_5,	ready_5_to_0;
wire    [`DATA_WIDTH-1:0]   data_5_to_10,	data_10_to_5;
wire                        valid_5_to_10,	valid_10_to_5;
wire                        ready_5_to_10,	ready_10_to_5;
wire    [`DATA_WIDTH-1:0]   data_10_to_15,	data_15_to_10;
wire                        valid_10_to_15,	valid_15_to_10;
wire                        ready_10_to_15,	ready_15_to_10;
wire    [`DATA_WIDTH-1:0]   data_15_to_20,	data_20_to_15;
wire                        valid_15_to_20,	valid_20_to_15;
wire                        ready_15_to_20,	ready_20_to_15;
wire    [`DATA_WIDTH-1:0]   data_1_to_6,	data_6_to_1;
wire                        valid_1_to_6,	valid_6_to_1;
wire                        ready_1_to_6,	ready_6_to_1;
wire    [`DATA_WIDTH-1:0]   data_6_to_11,	data_11_to_6;
wire                        valid_6_to_11,	valid_11_to_6;
wire                        ready_6_to_11,	ready_11_to_6;
wire    [`DATA_WIDTH-1:0]   data_11_to_16,	data_16_to_11;
wire                        valid_11_to_16,	valid_16_to_11;
wire                        ready_11_to_16,	ready_16_to_11;
wire    [`DATA_WIDTH-1:0]   data_16_to_21,	data_21_to_16;
wire                        valid_16_to_21,	valid_21_to_16;
wire                        ready_16_to_21,	ready_21_to_16;
wire    [`DATA_WIDTH-1:0]   data_2_to_7,	data_7_to_2;
wire                        valid_2_to_7,	valid_7_to_2;
wire                        ready_2_to_7,	ready_7_to_2;
wire    [`DATA_WIDTH-1:0]   data_7_to_12,	data_12_to_7;
wire                        valid_7_to_12,	valid_12_to_7;
wire                        ready_7_to_12,	ready_12_to_7;
wire    [`DATA_WIDTH-1:0]   data_12_to_17,	data_17_to_12;
wire                        valid_12_to_17,	valid_17_to_12;
wire                        ready_12_to_17,	ready_17_to_12;
wire    [`DATA_WIDTH-1:0]   data_17_to_22,	data_22_to_17;
wire                        valid_17_to_22,	valid_22_to_17;
wire                        ready_17_to_22,	ready_22_to_17;
wire    [`DATA_WIDTH-1:0]   data_3_to_8,	data_8_to_3;
wire                        valid_3_to_8,	valid_8_to_3;
wire                        ready_3_to_8,	ready_8_to_3;
wire    [`DATA_WIDTH-1:0]   data_8_to_13,	data_13_to_8;
wire                        valid_8_to_13,	valid_13_to_8;
wire                        ready_8_to_13,	ready_13_to_8;
wire    [`DATA_WIDTH-1:0]   data_13_to_18,	data_18_to_13;
wire                        valid_13_to_18,	valid_18_to_13;
wire                        ready_13_to_18,	ready_18_to_13;
wire    [`DATA_WIDTH-1:0]   data_18_to_23,	data_23_to_18;
wire                        valid_18_to_23,	valid_23_to_18;
wire                        ready_18_to_23,	ready_23_to_18;
wire    [`DATA_WIDTH-1:0]   data_4_to_9,	data_9_to_4;
wire                        valid_4_to_9,	valid_9_to_4;
wire                        ready_4_to_9,	ready_9_to_4;
wire    [`DATA_WIDTH-1:0]   data_9_to_14,	data_14_to_9;
wire                        valid_9_to_14,	valid_14_to_9;
wire                        ready_9_to_14,	ready_14_to_9;
wire    [`DATA_WIDTH-1:0]   data_14_to_19,	data_19_to_14;
wire                        valid_14_to_19,	valid_19_to_14;
wire                        ready_14_to_19,	ready_19_to_14;
wire    [`DATA_WIDTH-1:0]   data_19_to_24,	data_24_to_19;
wire                        valid_19_to_24,	valid_24_to_19;
wire                        ready_19_to_24,	ready_24_to_19;
    
router #(
    .ROUTER_ID_X        (0),
    .ROUTER_ID_Y        (0)
)router0(
    .CDCLK              (CDCLK),
    .CDRESETn           (CDRESETn),
    .CDIDATAW           (130'b0),
    .CDIVALIDW          (1'b0),
    .CDIREADYW          (),
    .CDODATAW           (),
    .CDOVALIDW          (),
    .CDOREADYW          (1'b0),
    .CDIDATAE           (data_1_to_0),
    .CDIVALIDE          (valid_1_to_0),
    .CDIREADYE          (ready_0_to_1),
    .CDODATAE           (data_0_to_1),
    .CDOVALIDE          (valid_0_to_1),
    .CDOREADYE          (ready_1_to_0),
    .CDIDATAL           (CDIDATA_X0_Y0),
    .CDIVALIDL          (CDIVALID_X0_Y0),
    .CDIREADYL          (CDIREADY_X0_Y0),
    .CDIDATAN           (130'b0),
    .CDIVALIDN          (1'b0),
    .CDIREADYN          (),
    .CDODATAN           (),
    .CDOVALIDN          (),
    .CDOREADYN          (1'b0),
    .CDIDATAS           (data_5_to_0),
    .CDIVALIDS          (valid_5_to_0),
    .CDIREADYS          (ready_0_to_5),
    .CDODATAS           (data_0_to_5),
    .CDOVALIDS          (valid_0_to_5),
    .CDOREADYS          (ready_5_to_0),
    .CDODATAL           (CDODATA_X0_Y0),
    .CDOVALIDL          (CDOVALID_X0_Y0),
    .CDOREADYL          (CDOREADY_X0_Y0)
);
    
router #(
    .ROUTER_ID_X        (0),
    .ROUTER_ID_Y        (1)
)router1(
    .CDCLK              (CDCLK),
    .CDRESETn           (CDRESETn),
    .CDIDATAW           (data_0_to_1),
    .CDIVALIDW          (valid_0_to_1),
    .CDIREADYW          (ready_1_to_0),
    .CDODATAW           (data_1_to_0),
    .CDOVALIDW          (valid_1_to_0),
    .CDOREADYW          (ready_0_to_1),
    .CDIDATAE           (data_2_to_1),
    .CDIVALIDE          (valid_2_to_1),
    .CDIREADYE          (ready_1_to_2),
    .CDODATAE           (data_1_to_2),
    .CDOVALIDE          (valid_1_to_2),
    .CDOREADYE          (ready_2_to_1),
    .CDIDATAL           (CDIDATA_X0_Y1),
    .CDIVALIDL          (CDIVALID_X0_Y1),
    .CDIREADYL          (CDIREADY_X0_Y1),
    .CDIDATAN           (130'b0),
    .CDIVALIDN          (1'b0),
    .CDIREADYN          (),
    .CDODATAN           (),
    .CDOVALIDN          (),
    .CDOREADYN          (1'b0),
    .CDIDATAS           (data_6_to_1),
    .CDIVALIDS          (valid_6_to_1),
    .CDIREADYS          (ready_1_to_6),
    .CDODATAS           (data_1_to_6),
    .CDOVALIDS          (valid_1_to_6),
    .CDOREADYS          (ready_6_to_1),
    .CDODATAL           (CDODATA_X0_Y1),
    .CDOVALIDL          (CDOVALID_X0_Y1),
    .CDOREADYL          (CDOREADY_X0_Y1)
);
    
router #(
    .ROUTER_ID_X        (0),
    .ROUTER_ID_Y        (2)
)router2(
    .CDCLK              (CDCLK),
    .CDRESETn           (CDRESETn),
    .CDIDATAW           (data_1_to_2),
    .CDIVALIDW          (valid_1_to_2),
    .CDIREADYW          (ready_2_to_1),
    .CDODATAW           (data_2_to_1),
    .CDOVALIDW          (valid_2_to_1),
    .CDOREADYW          (ready_1_to_2),
    .CDIDATAE           (data_3_to_2),
    .CDIVALIDE          (valid_3_to_2),
    .CDIREADYE          (ready_2_to_3),
    .CDODATAE           (data_2_to_3),
    .CDOVALIDE          (valid_2_to_3),
    .CDOREADYE          (ready_3_to_2),
    .CDIDATAL           (CDIDATA_X0_Y2),
    .CDIVALIDL          (CDIVALID_X0_Y2),
    .CDIREADYL          (CDIREADY_X0_Y2),
    .CDIDATAN           (130'b0),
    .CDIVALIDN          (1'b0),
    .CDIREADYN          (),
    .CDODATAN           (),
    .CDOVALIDN          (),
    .CDOREADYN          (1'b0),
    .CDIDATAS           (data_7_to_2),
    .CDIVALIDS          (valid_7_to_2),
    .CDIREADYS          (ready_2_to_7),
    .CDODATAS           (data_2_to_7),
    .CDOVALIDS          (valid_2_to_7),
    .CDOREADYS          (ready_7_to_2),
    .CDODATAL           (CDODATA_X0_Y2),
    .CDOVALIDL          (CDOVALID_X0_Y2),
    .CDOREADYL          (CDOREADY_X0_Y2)
);
    
router #(
    .ROUTER_ID_X        (0),
    .ROUTER_ID_Y        (3)
)router3(
    .CDCLK              (CDCLK),
    .CDRESETn           (CDRESETn),
    .CDIDATAW           (data_2_to_3),
    .CDIVALIDW          (valid_2_to_3),
    .CDIREADYW          (ready_3_to_2),
    .CDODATAW           (data_3_to_2),
    .CDOVALIDW          (valid_3_to_2),
    .CDOREADYW          (ready_2_to_3),
    .CDIDATAE           (data_4_to_3),
    .CDIVALIDE          (valid_4_to_3),
    .CDIREADYE          (ready_3_to_4),
    .CDODATAE           (data_3_to_4),
    .CDOVALIDE          (valid_3_to_4),
    .CDOREADYE          (ready_4_to_3),
    .CDIDATAL           (CDIDATA_X0_Y3),
    .CDIVALIDL          (CDIVALID_X0_Y3),
    .CDIREADYL          (CDIREADY_X0_Y3),
    .CDIDATAN           (130'b0),
    .CDIVALIDN          (1'b0),
    .CDIREADYN          (),
    .CDODATAN           (),
    .CDOVALIDN          (),
    .CDOREADYN          (1'b0),
    .CDIDATAS           (data_8_to_3),
    .CDIVALIDS          (valid_8_to_3),
    .CDIREADYS          (ready_3_to_8),
    .CDODATAS           (data_3_to_8),
    .CDOVALIDS          (valid_3_to_8),
    .CDOREADYS          (ready_8_to_3),
    .CDODATAL           (CDODATA_X0_Y3),
    .CDOVALIDL          (CDOVALID_X0_Y3),
    .CDOREADYL          (CDOREADY_X0_Y3)
);
    
router #(
    .ROUTER_ID_X        (0),
    .ROUTER_ID_Y        (4)
)router4(
    .CDCLK              (CDCLK),
    .CDRESETn           (CDRESETn),
    .CDIDATAW           (data_3_to_4),
    .CDIVALIDW          (valid_3_to_4),
    .CDIREADYW          (ready_4_to_3),
    .CDODATAW           (data_4_to_3),
    .CDOVALIDW          (valid_4_to_3),
    .CDOREADYW          (ready_3_to_4),
    .CDIDATAE           (130'b0),
    .CDIVALIDE          (1'b0),
    .CDIREADYE          (),
    .CDODATAE           (),
    .CDOVALIDE          (),
    .CDOREADYE          (1'b0),
    .CDIDATAL           (CDIDATA_X0_Y4),
    .CDIVALIDL          (CDIVALID_X0_Y4),
    .CDIREADYL          (CDIREADY_X0_Y4),
    .CDIDATAN           (130'b0),
    .CDIVALIDN          (1'b0),
    .CDIREADYN          (),
    .CDODATAN           (),
    .CDOVALIDN          (),
    .CDOREADYN          (1'b0),
    .CDIDATAS           (data_9_to_4),
    .CDIVALIDS          (valid_9_to_4),
    .CDIREADYS          (ready_4_to_9),
    .CDODATAS           (data_4_to_9),
    .CDOVALIDS          (valid_4_to_9),
    .CDOREADYS          (ready_9_to_4),
    .CDODATAL           (CDODATA_X0_Y4),
    .CDOVALIDL          (CDOVALID_X0_Y4),
    .CDOREADYL          (CDOREADY_X0_Y4)
);
    
router #(
    .ROUTER_ID_X        (1),
    .ROUTER_ID_Y        (0)
)router5(
    .CDCLK              (CDCLK),
    .CDRESETn           (CDRESETn),
    .CDIDATAW           (130'b0),
    .CDIVALIDW          (1'b0),
    .CDIREADYW          (),
    .CDODATAW           (),
    .CDOVALIDW          (),
    .CDOREADYW          (1'b0),
    .CDIDATAE           (data_6_to_5),
    .CDIVALIDE          (valid_6_to_5),
    .CDIREADYE          (ready_5_to_6),
    .CDODATAE           (data_5_to_6),
    .CDOVALIDE          (valid_5_to_6),
    .CDOREADYE          (ready_6_to_5),
    .CDIDATAL           (CDIDATA_X1_Y0),
    .CDIVALIDL          (CDIVALID_X1_Y0),
    .CDIREADYL          (CDIREADY_X1_Y0),
    .CDIDATAN           (data_0_to_5),
    .CDIVALIDN          (valid_0_to_5),
    .CDIREADYN          (ready_5_to_0),
    .CDODATAN           (data_5_to_0),
    .CDOVALIDN          (valid_5_to_0),
    .CDOREADYN          (ready_0_to_5),
    .CDIDATAS           (data_10_to_5),
    .CDIVALIDS          (valid_10_to_5),
    .CDIREADYS          (ready_5_to_10),
    .CDODATAS           (data_5_to_10),
    .CDOVALIDS          (valid_5_to_10),
    .CDOREADYS          (ready_10_to_5),
    .CDODATAL           (CDODATA_X1_Y0),
    .CDOVALIDL          (CDOVALID_X1_Y0),
    .CDOREADYL          (CDOREADY_X1_Y0)
);
    
router #(
    .ROUTER_ID_X        (1),
    .ROUTER_ID_Y        (1)
)router6(
    .CDCLK              (CDCLK),
    .CDRESETn           (CDRESETn),
    .CDIDATAW           (data_5_to_6),
    .CDIVALIDW          (valid_5_to_6),
    .CDIREADYW          (ready_6_to_5),
    .CDODATAW           (data_6_to_5),
    .CDOVALIDW          (valid_6_to_5),
    .CDOREADYW          (ready_5_to_6),
    .CDIDATAE           (data_7_to_6),
    .CDIVALIDE          (valid_7_to_6),
    .CDIREADYE          (ready_6_to_7),
    .CDODATAE           (data_6_to_7),
    .CDOVALIDE          (valid_6_to_7),
    .CDOREADYE          (ready_7_to_6),
    .CDIDATAL           (CDIDATA_X1_Y1),
    .CDIVALIDL          (CDIVALID_X1_Y1),
    .CDIREADYL          (CDIREADY_X1_Y1),
    .CDIDATAN           (data_1_to_6),
    .CDIVALIDN          (valid_1_to_6),
    .CDIREADYN          (ready_6_to_1),
    .CDODATAN           (data_6_to_1),
    .CDOVALIDN          (valid_6_to_1),
    .CDOREADYN          (ready_1_to_6),
    .CDIDATAS           (data_11_to_6),
    .CDIVALIDS          (valid_11_to_6),
    .CDIREADYS          (ready_6_to_11),
    .CDODATAS           (data_6_to_11),
    .CDOVALIDS          (valid_6_to_11),
    .CDOREADYS          (ready_11_to_6),
    .CDODATAL           (CDODATA_X1_Y1),
    .CDOVALIDL          (CDOVALID_X1_Y1),
    .CDOREADYL          (CDOREADY_X1_Y1)
);
    
router #(
    .ROUTER_ID_X        (1),
    .ROUTER_ID_Y        (2)
)router7(
    .CDCLK              (CDCLK),
    .CDRESETn           (CDRESETn),
    .CDIDATAW           (data_6_to_7),
    .CDIVALIDW          (valid_6_to_7),
    .CDIREADYW          (ready_7_to_6),
    .CDODATAW           (data_7_to_6),
    .CDOVALIDW          (valid_7_to_6),
    .CDOREADYW          (ready_6_to_7),
    .CDIDATAE           (data_8_to_7),
    .CDIVALIDE          (valid_8_to_7),
    .CDIREADYE          (ready_7_to_8),
    .CDODATAE           (data_7_to_8),
    .CDOVALIDE          (valid_7_to_8),
    .CDOREADYE          (ready_8_to_7),
    .CDIDATAL           (CDIDATA_X1_Y2),
    .CDIVALIDL          (CDIVALID_X1_Y2),
    .CDIREADYL          (CDIREADY_X1_Y2),
    .CDIDATAN           (data_2_to_7),
    .CDIVALIDN          (valid_2_to_7),
    .CDIREADYN          (ready_7_to_2),
    .CDODATAN           (data_7_to_2),
    .CDOVALIDN          (valid_7_to_2),
    .CDOREADYN          (ready_2_to_7),
    .CDIDATAS           (data_12_to_7),
    .CDIVALIDS          (valid_12_to_7),
    .CDIREADYS          (ready_7_to_12),
    .CDODATAS           (data_7_to_12),
    .CDOVALIDS          (valid_7_to_12),
    .CDOREADYS          (ready_12_to_7),
    .CDODATAL           (CDODATA_X1_Y2),
    .CDOVALIDL          (CDOVALID_X1_Y2),
    .CDOREADYL          (CDOREADY_X1_Y2)
);
    
router #(
    .ROUTER_ID_X        (1),
    .ROUTER_ID_Y        (3)
)router8(
    .CDCLK              (CDCLK),
    .CDRESETn           (CDRESETn),
    .CDIDATAW           (data_7_to_8),
    .CDIVALIDW          (valid_7_to_8),
    .CDIREADYW          (ready_8_to_7),
    .CDODATAW           (data_8_to_7),
    .CDOVALIDW          (valid_8_to_7),
    .CDOREADYW          (ready_7_to_8),
    .CDIDATAE           (data_9_to_8),
    .CDIVALIDE          (valid_9_to_8),
    .CDIREADYE          (ready_8_to_9),
    .CDODATAE           (data_8_to_9),
    .CDOVALIDE          (valid_8_to_9),
    .CDOREADYE          (ready_9_to_8),
    .CDIDATAL           (CDIDATA_X1_Y3),
    .CDIVALIDL          (CDIVALID_X1_Y3),
    .CDIREADYL          (CDIREADY_X1_Y3),
    .CDIDATAN           (data_3_to_8),
    .CDIVALIDN          (valid_3_to_8),
    .CDIREADYN          (ready_8_to_3),
    .CDODATAN           (data_8_to_3),
    .CDOVALIDN          (valid_8_to_3),
    .CDOREADYN          (ready_3_to_8),
    .CDIDATAS           (data_13_to_8),
    .CDIVALIDS          (valid_13_to_8),
    .CDIREADYS          (ready_8_to_13),
    .CDODATAS           (data_8_to_13),
    .CDOVALIDS          (valid_8_to_13),
    .CDOREADYS          (ready_13_to_8),
    .CDODATAL           (CDODATA_X1_Y3),
    .CDOVALIDL          (CDOVALID_X1_Y3),
    .CDOREADYL          (CDOREADY_X1_Y3)
);
    
router #(
    .ROUTER_ID_X        (1),
    .ROUTER_ID_Y        (4)
)router9(
    .CDCLK              (CDCLK),
    .CDRESETn           (CDRESETn),
    .CDIDATAW           (data_8_to_9),
    .CDIVALIDW          (valid_8_to_9),
    .CDIREADYW          (ready_9_to_8),
    .CDODATAW           (data_9_to_8),
    .CDOVALIDW          (valid_9_to_8),
    .CDOREADYW          (ready_8_to_9),
    .CDIDATAE           (130'b0),
    .CDIVALIDE          (1'b0),
    .CDIREADYE          (),
    .CDODATAE           (),
    .CDOVALIDE          (),
    .CDOREADYE          (1'b0),
    .CDIDATAL           (CDIDATA_X1_Y4),
    .CDIVALIDL          (CDIVALID_X1_Y4),
    .CDIREADYL          (CDIREADY_X1_Y4),
    .CDIDATAN           (data_4_to_9),
    .CDIVALIDN          (valid_4_to_9),
    .CDIREADYN          (ready_9_to_4),
    .CDODATAN           (data_9_to_4),
    .CDOVALIDN          (valid_9_to_4),
    .CDOREADYN          (ready_4_to_9),
    .CDIDATAS           (data_14_to_9),
    .CDIVALIDS          (valid_14_to_9),
    .CDIREADYS          (ready_9_to_14),
    .CDODATAS           (data_9_to_14),
    .CDOVALIDS          (valid_9_to_14),
    .CDOREADYS          (ready_14_to_9),
    .CDODATAL           (CDODATA_X1_Y4),
    .CDOVALIDL          (CDOVALID_X1_Y4),
    .CDOREADYL          (CDOREADY_X1_Y4)
);
    
router #(
    .ROUTER_ID_X        (2),
    .ROUTER_ID_Y        (0)
)router10(
    .CDCLK              (CDCLK),
    .CDRESETn           (CDRESETn),
    .CDIDATAW           (130'b0),
    .CDIVALIDW          (1'b0),
    .CDIREADYW          (),
    .CDODATAW           (),
    .CDOVALIDW          (),
    .CDOREADYW          (1'b0),
    .CDIDATAE           (data_11_to_10),
    .CDIVALIDE          (valid_11_to_10),
    .CDIREADYE          (ready_10_to_11),
    .CDODATAE           (data_10_to_11),
    .CDOVALIDE          (valid_10_to_11),
    .CDOREADYE          (ready_11_to_10),
    .CDIDATAL           (CDIDATA_X2_Y0),
    .CDIVALIDL          (CDIVALID_X2_Y0),
    .CDIREADYL          (CDIREADY_X2_Y0),
    .CDIDATAN           (data_5_to_10),
    .CDIVALIDN          (valid_5_to_10),
    .CDIREADYN          (ready_10_to_5),
    .CDODATAN           (data_10_to_5),
    .CDOVALIDN          (valid_10_to_5),
    .CDOREADYN          (ready_5_to_10),
    .CDIDATAS           (data_15_to_10),
    .CDIVALIDS          (valid_15_to_10),
    .CDIREADYS          (ready_10_to_15),
    .CDODATAS           (data_10_to_15),
    .CDOVALIDS          (valid_10_to_15),
    .CDOREADYS          (ready_15_to_10),
    .CDODATAL           (CDODATA_X2_Y0),
    .CDOVALIDL          (CDOVALID_X2_Y0),
    .CDOREADYL          (CDOREADY_X2_Y0)
);
    
router #(
    .ROUTER_ID_X        (2),
    .ROUTER_ID_Y        (1)
)router11(
    .CDCLK              (CDCLK),
    .CDRESETn           (CDRESETn),
    .CDIDATAW           (data_10_to_11),
    .CDIVALIDW          (valid_10_to_11),
    .CDIREADYW          (ready_11_to_10),
    .CDODATAW           (data_11_to_10),
    .CDOVALIDW          (valid_11_to_10),
    .CDOREADYW          (ready_10_to_11),
    .CDIDATAE           (data_12_to_11),
    .CDIVALIDE          (valid_12_to_11),
    .CDIREADYE          (ready_11_to_12),
    .CDODATAE           (data_11_to_12),
    .CDOVALIDE          (valid_11_to_12),
    .CDOREADYE          (ready_12_to_11),
    .CDIDATAL           (CDIDATA_X2_Y1),
    .CDIVALIDL          (CDIVALID_X2_Y1),
    .CDIREADYL          (CDIREADY_X2_Y1),
    .CDIDATAN           (data_6_to_11),
    .CDIVALIDN          (valid_6_to_11),
    .CDIREADYN          (ready_11_to_6),
    .CDODATAN           (data_11_to_6),
    .CDOVALIDN          (valid_11_to_6),
    .CDOREADYN          (ready_6_to_11),
    .CDIDATAS           (data_16_to_11),
    .CDIVALIDS          (valid_16_to_11),
    .CDIREADYS          (ready_11_to_16),
    .CDODATAS           (data_11_to_16),
    .CDOVALIDS          (valid_11_to_16),
    .CDOREADYS          (ready_16_to_11),
    .CDODATAL           (CDODATA_X2_Y1),
    .CDOVALIDL          (CDOVALID_X2_Y1),
    .CDOREADYL          (CDOREADY_X2_Y1)
);
    
router #(
    .ROUTER_ID_X        (2),
    .ROUTER_ID_Y        (2)
)router12(
    .CDCLK              (CDCLK),
    .CDRESETn           (CDRESETn),
    .CDIDATAW           (data_11_to_12),
    .CDIVALIDW          (valid_11_to_12),
    .CDIREADYW          (ready_12_to_11),
    .CDODATAW           (data_12_to_11),
    .CDOVALIDW          (valid_12_to_11),
    .CDOREADYW          (ready_11_to_12),
    .CDIDATAE           (data_13_to_12),
    .CDIVALIDE          (valid_13_to_12),
    .CDIREADYE          (ready_12_to_13),
    .CDODATAE           (data_12_to_13),
    .CDOVALIDE          (valid_12_to_13),
    .CDOREADYE          (ready_13_to_12),
    .CDIDATAL           (CDIDATA_X2_Y2),
    .CDIVALIDL          (CDIVALID_X2_Y2),
    .CDIREADYL          (CDIREADY_X2_Y2),
    .CDIDATAN           (data_7_to_12),
    .CDIVALIDN          (valid_7_to_12),
    .CDIREADYN          (ready_12_to_7),
    .CDODATAN           (data_12_to_7),
    .CDOVALIDN          (valid_12_to_7),
    .CDOREADYN          (ready_7_to_12),
    .CDIDATAS           (data_17_to_12),
    .CDIVALIDS          (valid_17_to_12),
    .CDIREADYS          (ready_12_to_17),
    .CDODATAS           (data_12_to_17),
    .CDOVALIDS          (valid_12_to_17),
    .CDOREADYS          (ready_17_to_12),
    .CDODATAL           (CDODATA_X2_Y2),
    .CDOVALIDL          (CDOVALID_X2_Y2),
    .CDOREADYL          (CDOREADY_X2_Y2)
);
    
router #(
    .ROUTER_ID_X        (2),
    .ROUTER_ID_Y        (3)
)router13(
    .CDCLK              (CDCLK),
    .CDRESETn           (CDRESETn),
    .CDIDATAW           (data_12_to_13),
    .CDIVALIDW          (valid_12_to_13),
    .CDIREADYW          (ready_13_to_12),
    .CDODATAW           (data_13_to_12),
    .CDOVALIDW          (valid_13_to_12),
    .CDOREADYW          (ready_12_to_13),
    .CDIDATAE           (data_14_to_13),
    .CDIVALIDE          (valid_14_to_13),
    .CDIREADYE          (ready_13_to_14),
    .CDODATAE           (data_13_to_14),
    .CDOVALIDE          (valid_13_to_14),
    .CDOREADYE          (ready_14_to_13),
    .CDIDATAL           (CDIDATA_X2_Y3),
    .CDIVALIDL          (CDIVALID_X2_Y3),
    .CDIREADYL          (CDIREADY_X2_Y3),
    .CDIDATAN           (data_8_to_13),
    .CDIVALIDN          (valid_8_to_13),
    .CDIREADYN          (ready_13_to_8),
    .CDODATAN           (data_13_to_8),
    .CDOVALIDN          (valid_13_to_8),
    .CDOREADYN          (ready_8_to_13),
    .CDIDATAS           (data_18_to_13),
    .CDIVALIDS          (valid_18_to_13),
    .CDIREADYS          (ready_13_to_18),
    .CDODATAS           (data_13_to_18),
    .CDOVALIDS          (valid_13_to_18),
    .CDOREADYS          (ready_18_to_13),
    .CDODATAL           (CDODATA_X2_Y3),
    .CDOVALIDL          (CDOVALID_X2_Y3),
    .CDOREADYL          (CDOREADY_X2_Y3)
);
    
router #(
    .ROUTER_ID_X        (2),
    .ROUTER_ID_Y        (4)
)router14(
    .CDCLK              (CDCLK),
    .CDRESETn           (CDRESETn),
    .CDIDATAW           (data_13_to_14),
    .CDIVALIDW          (valid_13_to_14),
    .CDIREADYW          (ready_14_to_13),
    .CDODATAW           (data_14_to_13),
    .CDOVALIDW          (valid_14_to_13),
    .CDOREADYW          (ready_13_to_14),
    .CDIDATAE           (130'b0),
    .CDIVALIDE          (1'b0),
    .CDIREADYE          (),
    .CDODATAE           (),
    .CDOVALIDE          (),
    .CDOREADYE          (1'b0),
    .CDIDATAL           (CDIDATA_X2_Y4),
    .CDIVALIDL          (CDIVALID_X2_Y4),
    .CDIREADYL          (CDIREADY_X2_Y4),
    .CDIDATAN           (data_9_to_14),
    .CDIVALIDN          (valid_9_to_14),
    .CDIREADYN          (ready_14_to_9),
    .CDODATAN           (data_14_to_9),
    .CDOVALIDN          (valid_14_to_9),
    .CDOREADYN          (ready_9_to_14),
    .CDIDATAS           (data_19_to_14),
    .CDIVALIDS          (valid_19_to_14),
    .CDIREADYS          (ready_14_to_19),
    .CDODATAS           (data_14_to_19),
    .CDOVALIDS          (valid_14_to_19),
    .CDOREADYS          (ready_19_to_14),
    .CDODATAL           (CDODATA_X2_Y4),
    .CDOVALIDL          (CDOVALID_X2_Y4),
    .CDOREADYL          (CDOREADY_X2_Y4)
);
    
router #(
    .ROUTER_ID_X        (3),
    .ROUTER_ID_Y        (0)
)router15(
    .CDCLK              (CDCLK),
    .CDRESETn           (CDRESETn),
    .CDIDATAW           (130'b0),
    .CDIVALIDW          (1'b0),
    .CDIREADYW          (),
    .CDODATAW           (),
    .CDOVALIDW          (),
    .CDOREADYW          (1'b0),
    .CDIDATAE           (data_16_to_15),
    .CDIVALIDE          (valid_16_to_15),
    .CDIREADYE          (ready_15_to_16),
    .CDODATAE           (data_15_to_16),
    .CDOVALIDE          (valid_15_to_16),
    .CDOREADYE          (ready_16_to_15),
    .CDIDATAL           (CDIDATA_X3_Y0),
    .CDIVALIDL          (CDIVALID_X3_Y0),
    .CDIREADYL          (CDIREADY_X3_Y0),
    .CDIDATAN           (data_10_to_15),
    .CDIVALIDN          (valid_10_to_15),
    .CDIREADYN          (ready_15_to_10),
    .CDODATAN           (data_15_to_10),
    .CDOVALIDN          (valid_15_to_10),
    .CDOREADYN          (ready_10_to_15),
    .CDIDATAS           (data_20_to_15),
    .CDIVALIDS          (valid_20_to_15),
    .CDIREADYS          (ready_15_to_20),
    .CDODATAS           (data_15_to_20),
    .CDOVALIDS          (valid_15_to_20),
    .CDOREADYS          (ready_20_to_15),
    .CDODATAL           (CDODATA_X3_Y0),
    .CDOVALIDL          (CDOVALID_X3_Y0),
    .CDOREADYL          (CDOREADY_X3_Y0)
);
    
router #(
    .ROUTER_ID_X        (3),
    .ROUTER_ID_Y        (1)
)router16(
    .CDCLK              (CDCLK),
    .CDRESETn           (CDRESETn),
    .CDIDATAW           (data_15_to_16),
    .CDIVALIDW          (valid_15_to_16),
    .CDIREADYW          (ready_16_to_15),
    .CDODATAW           (data_16_to_15),
    .CDOVALIDW          (valid_16_to_15),
    .CDOREADYW          (ready_15_to_16),
    .CDIDATAE           (data_17_to_16),
    .CDIVALIDE          (valid_17_to_16),
    .CDIREADYE          (ready_16_to_17),
    .CDODATAE           (data_16_to_17),
    .CDOVALIDE          (valid_16_to_17),
    .CDOREADYE          (ready_17_to_16),
    .CDIDATAL           (CDIDATA_X3_Y1),
    .CDIVALIDL          (CDIVALID_X3_Y1),
    .CDIREADYL          (CDIREADY_X3_Y1),
    .CDIDATAN           (data_11_to_16),
    .CDIVALIDN          (valid_11_to_16),
    .CDIREADYN          (ready_16_to_11),
    .CDODATAN           (data_16_to_11),
    .CDOVALIDN          (valid_16_to_11),
    .CDOREADYN          (ready_11_to_16),
    .CDIDATAS           (data_21_to_16),
    .CDIVALIDS          (valid_21_to_16),
    .CDIREADYS          (ready_16_to_21),
    .CDODATAS           (data_16_to_21),
    .CDOVALIDS          (valid_16_to_21),
    .CDOREADYS          (ready_21_to_16),
    .CDODATAL           (CDODATA_X3_Y1),
    .CDOVALIDL          (CDOVALID_X3_Y1),
    .CDOREADYL          (CDOREADY_X3_Y1)
);
    
router #(
    .ROUTER_ID_X        (3),
    .ROUTER_ID_Y        (2)
)router17(
    .CDCLK              (CDCLK),
    .CDRESETn           (CDRESETn),
    .CDIDATAW           (data_16_to_17),
    .CDIVALIDW          (valid_16_to_17),
    .CDIREADYW          (ready_17_to_16),
    .CDODATAW           (data_17_to_16),
    .CDOVALIDW          (valid_17_to_16),
    .CDOREADYW          (ready_16_to_17),
    .CDIDATAE           (data_18_to_17),
    .CDIVALIDE          (valid_18_to_17),
    .CDIREADYE          (ready_17_to_18),
    .CDODATAE           (data_17_to_18),
    .CDOVALIDE          (valid_17_to_18),
    .CDOREADYE          (ready_18_to_17),
    .CDIDATAL           (CDIDATA_X3_Y2),
    .CDIVALIDL          (CDIVALID_X3_Y2),
    .CDIREADYL          (CDIREADY_X3_Y2),
    .CDIDATAN           (data_12_to_17),
    .CDIVALIDN          (valid_12_to_17),
    .CDIREADYN          (ready_17_to_12),
    .CDODATAN           (data_17_to_12),
    .CDOVALIDN          (valid_17_to_12),
    .CDOREADYN          (ready_12_to_17),
    .CDIDATAS           (data_22_to_17),
    .CDIVALIDS          (valid_22_to_17),
    .CDIREADYS          (ready_17_to_22),
    .CDODATAS           (data_17_to_22),
    .CDOVALIDS          (valid_17_to_22),
    .CDOREADYS          (ready_22_to_17),
    .CDODATAL           (CDODATA_X3_Y2),
    .CDOVALIDL          (CDOVALID_X3_Y2),
    .CDOREADYL          (CDOREADY_X3_Y2)
);
    
router #(
    .ROUTER_ID_X        (3),
    .ROUTER_ID_Y        (3)
)router18(
    .CDCLK              (CDCLK),
    .CDRESETn           (CDRESETn),
    .CDIDATAW           (data_17_to_18),
    .CDIVALIDW          (valid_17_to_18),
    .CDIREADYW          (ready_18_to_17),
    .CDODATAW           (data_18_to_17),
    .CDOVALIDW          (valid_18_to_17),
    .CDOREADYW          (ready_17_to_18),
    .CDIDATAE           (data_19_to_18),
    .CDIVALIDE          (valid_19_to_18),
    .CDIREADYE          (ready_18_to_19),
    .CDODATAE           (data_18_to_19),
    .CDOVALIDE          (valid_18_to_19),
    .CDOREADYE          (ready_19_to_18),
    .CDIDATAL           (CDIDATA_X3_Y3),
    .CDIVALIDL          (CDIVALID_X3_Y3),
    .CDIREADYL          (CDIREADY_X3_Y3),
    .CDIDATAN           (data_13_to_18),
    .CDIVALIDN          (valid_13_to_18),
    .CDIREADYN          (ready_18_to_13),
    .CDODATAN           (data_18_to_13),
    .CDOVALIDN          (valid_18_to_13),
    .CDOREADYN          (ready_13_to_18),
    .CDIDATAS           (data_23_to_18),
    .CDIVALIDS          (valid_23_to_18),
    .CDIREADYS          (ready_18_to_23),
    .CDODATAS           (data_18_to_23),
    .CDOVALIDS          (valid_18_to_23),
    .CDOREADYS          (ready_23_to_18),
    .CDODATAL           (CDODATA_X3_Y3),
    .CDOVALIDL          (CDOVALID_X3_Y3),
    .CDOREADYL          (CDOREADY_X3_Y3)
);
    
router #(
    .ROUTER_ID_X        (3),
    .ROUTER_ID_Y        (4)
)router19(
    .CDCLK              (CDCLK),
    .CDRESETn           (CDRESETn),
    .CDIDATAW           (data_18_to_19),
    .CDIVALIDW          (valid_18_to_19),
    .CDIREADYW          (ready_19_to_18),
    .CDODATAW           (data_19_to_18),
    .CDOVALIDW          (valid_19_to_18),
    .CDOREADYW          (ready_18_to_19),
    .CDIDATAE           (130'b0),
    .CDIVALIDE          (1'b0),
    .CDIREADYE          (),
    .CDODATAE           (),
    .CDOVALIDE          (),
    .CDOREADYE          (1'b0),
    .CDIDATAL           (CDIDATA_X3_Y4),
    .CDIVALIDL          (CDIVALID_X3_Y4),
    .CDIREADYL          (CDIREADY_X3_Y4),
    .CDIDATAN           (data_14_to_19),
    .CDIVALIDN          (valid_14_to_19),
    .CDIREADYN          (ready_19_to_14),
    .CDODATAN           (data_19_to_14),
    .CDOVALIDN          (valid_19_to_14),
    .CDOREADYN          (ready_14_to_19),
    .CDIDATAS           (data_24_to_19),
    .CDIVALIDS          (valid_24_to_19),
    .CDIREADYS          (ready_19_to_24),
    .CDODATAS           (data_19_to_24),
    .CDOVALIDS          (valid_19_to_24),
    .CDOREADYS          (ready_24_to_19),
    .CDODATAL           (CDODATA_X3_Y4),
    .CDOVALIDL          (CDOVALID_X3_Y4),
    .CDOREADYL          (CDOREADY_X3_Y4)
);
    
router #(
    .ROUTER_ID_X        (4),
    .ROUTER_ID_Y        (0)
)router20(
    .CDCLK              (CDCLK),
    .CDRESETn           (CDRESETn),
    .CDIDATAW           (130'b0),
    .CDIVALIDW          (1'b0),
    .CDIREADYW          (),
    .CDODATAW           (),
    .CDOVALIDW          (),
    .CDOREADYW          (1'b0),
    .CDIDATAE           (data_21_to_20),
    .CDIVALIDE          (valid_21_to_20),
    .CDIREADYE          (ready_20_to_21),
    .CDODATAE           (data_20_to_21),
    .CDOVALIDE          (valid_20_to_21),
    .CDOREADYE          (ready_21_to_20),
    .CDIDATAL           (CDIDATA_X4_Y0),
    .CDIVALIDL          (CDIVALID_X4_Y0),
    .CDIREADYL          (CDIREADY_X4_Y0),
    .CDIDATAN           (data_15_to_20),
    .CDIVALIDN          (valid_15_to_20),
    .CDIREADYN          (ready_20_to_15),
    .CDODATAN           (data_20_to_15),
    .CDOVALIDN          (valid_20_to_15),
    .CDOREADYN          (ready_15_to_20),
    .CDIDATAS           (130'b0),
    .CDIVALIDS          (1'b0),
    .CDIREADYS          (),
    .CDODATAS           (),
    .CDOVALIDS          (),
    .CDOREADYS          (1'b0),
    .CDODATAL           (CDODATA_X4_Y0),
    .CDOVALIDL          (CDOVALID_X4_Y0),
    .CDOREADYL          (CDOREADY_X4_Y0)
);
    
router #(
    .ROUTER_ID_X        (4),
    .ROUTER_ID_Y        (1)
)router21(
    .CDCLK              (CDCLK),
    .CDRESETn           (CDRESETn),
    .CDIDATAW           (data_20_to_21),
    .CDIVALIDW          (valid_20_to_21),
    .CDIREADYW          (ready_21_to_20),
    .CDODATAW           (data_21_to_20),
    .CDOVALIDW          (valid_21_to_20),
    .CDOREADYW          (ready_20_to_21),
    .CDIDATAE           (data_22_to_21),
    .CDIVALIDE          (valid_22_to_21),
    .CDIREADYE          (ready_21_to_22),
    .CDODATAE           (data_21_to_22),
    .CDOVALIDE          (valid_21_to_22),
    .CDOREADYE          (ready_22_to_21),
    .CDIDATAL           (CDIDATA_X4_Y1),
    .CDIVALIDL          (CDIVALID_X4_Y1),
    .CDIREADYL          (CDIREADY_X4_Y1),
    .CDIDATAN           (data_16_to_21),
    .CDIVALIDN          (valid_16_to_21),
    .CDIREADYN          (ready_21_to_16),
    .CDODATAN           (data_21_to_16),
    .CDOVALIDN          (valid_21_to_16),
    .CDOREADYN          (ready_16_to_21),
    .CDIDATAS           (130'b0),
    .CDIVALIDS          (1'b0),
    .CDIREADYS          (),
    .CDODATAS           (),
    .CDOVALIDS          (),
    .CDOREADYS          (1'b0),
    .CDODATAL           (CDODATA_X4_Y1),
    .CDOVALIDL          (CDOVALID_X4_Y1),
    .CDOREADYL          (CDOREADY_X4_Y1)
);
    
router #(
    .ROUTER_ID_X        (4),
    .ROUTER_ID_Y        (2)
)router22(
    .CDCLK              (CDCLK),
    .CDRESETn           (CDRESETn),
    .CDIDATAW           (data_21_to_22),
    .CDIVALIDW          (valid_21_to_22),
    .CDIREADYW          (ready_22_to_21),
    .CDODATAW           (data_22_to_21),
    .CDOVALIDW          (valid_22_to_21),
    .CDOREADYW          (ready_21_to_22),
    .CDIDATAE           (data_23_to_22),
    .CDIVALIDE          (valid_23_to_22),
    .CDIREADYE          (ready_22_to_23),
    .CDODATAE           (data_22_to_23),
    .CDOVALIDE          (valid_22_to_23),
    .CDOREADYE          (ready_23_to_22),
    .CDIDATAL           (CDIDATA_X4_Y2),
    .CDIVALIDL          (CDIVALID_X4_Y2),
    .CDIREADYL          (CDIREADY_X4_Y2),
    .CDIDATAN           (data_17_to_22),
    .CDIVALIDN          (valid_17_to_22),
    .CDIREADYN          (ready_22_to_17),
    .CDODATAN           (data_22_to_17),
    .CDOVALIDN          (valid_22_to_17),
    .CDOREADYN          (ready_17_to_22),
    .CDIDATAS           (130'b0),
    .CDIVALIDS          (1'b0),
    .CDIREADYS          (),
    .CDODATAS           (),
    .CDOVALIDS          (),
    .CDOREADYS          (1'b0),
    .CDODATAL           (CDODATA_X4_Y2),
    .CDOVALIDL          (CDOVALID_X4_Y2),
    .CDOREADYL          (CDOREADY_X4_Y2)
);
    
router #(
    .ROUTER_ID_X        (4),
    .ROUTER_ID_Y        (3)
)router23(
    .CDCLK              (CDCLK),
    .CDRESETn           (CDRESETn),
    .CDIDATAW           (data_22_to_23),
    .CDIVALIDW          (valid_22_to_23),
    .CDIREADYW          (ready_23_to_22),
    .CDODATAW           (data_23_to_22),
    .CDOVALIDW          (valid_23_to_22),
    .CDOREADYW          (ready_22_to_23),
    .CDIDATAE           (data_24_to_23),
    .CDIVALIDE          (valid_24_to_23),
    .CDIREADYE          (ready_23_to_24),
    .CDODATAE           (data_23_to_24),
    .CDOVALIDE          (valid_23_to_24),
    .CDOREADYE          (ready_24_to_23),
    .CDIDATAL           (CDIDATA_X4_Y3),
    .CDIVALIDL          (CDIVALID_X4_Y3),
    .CDIREADYL          (CDIREADY_X4_Y3),
    .CDIDATAN           (data_18_to_23),
    .CDIVALIDN          (valid_18_to_23),
    .CDIREADYN          (ready_23_to_18),
    .CDODATAN           (data_23_to_18),
    .CDOVALIDN          (valid_23_to_18),
    .CDOREADYN          (ready_18_to_23),
    .CDIDATAS           (130'b0),
    .CDIVALIDS          (1'b0),
    .CDIREADYS          (),
    .CDODATAS           (),
    .CDOVALIDS          (),
    .CDOREADYS          (1'b0),
    .CDODATAL           (CDODATA_X4_Y3),
    .CDOVALIDL          (CDOVALID_X4_Y3),
    .CDOREADYL          (CDOREADY_X4_Y3)
);
    
router #(
    .ROUTER_ID_X        (4),
    .ROUTER_ID_Y        (4)
)router24(
    .CDCLK              (CDCLK),
    .CDRESETn           (CDRESETn),
    .CDIDATAW           (data_23_to_24),
    .CDIVALIDW          (valid_23_to_24),
    .CDIREADYW          (ready_24_to_23),
    .CDODATAW           (data_24_to_23),
    .CDOVALIDW          (valid_24_to_23),
    .CDOREADYW          (ready_23_to_24),
    .CDIDATAE           (130'b0),
    .CDIVALIDE          (1'b0),
    .CDIREADYE          (),
    .CDODATAE           (),
    .CDOVALIDE          (),
    .CDOREADYE          (1'b0),
    .CDIDATAL           (CDIDATA_X4_Y4),
    .CDIVALIDL          (CDIVALID_X4_Y4),
    .CDIREADYL          (CDIREADY_X4_Y4),
    .CDIDATAN           (data_19_to_24),
    .CDIVALIDN          (valid_19_to_24),
    .CDIREADYN          (ready_24_to_19),
    .CDODATAN           (data_24_to_19),
    .CDOVALIDN          (valid_24_to_19),
    .CDOREADYN          (ready_19_to_24),
    .CDIDATAS           (130'b0),
    .CDIVALIDS          (1'b0),
    .CDIREADYS          (),
    .CDODATAS           (),
    .CDOVALIDS          (),
    .CDOREADYS          (1'b0),
    .CDODATAL           (CDODATA_X4_Y4),
    .CDOVALIDL          (CDOVALID_X4_Y4),
    .CDOREADYL          (CDOREADY_X4_Y4)
);

endmodule
