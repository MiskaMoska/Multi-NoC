`include "param.vh"

module NoP(
    input       wire                                CDCLK,
    input       wire                                CPCLK,
    input       wire                                CDRESETn,
    
    //==============================================================//
    //                                                              /
    //                           NoD0                               /
    //                                                              /
    //==============================================================//
    //router0
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X0_Y0_D0,
    input       wire                                CDIVALID_X0_Y0_D0,
    output      wire                                CDIREADY_X0_Y0_D0,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X0_Y0_D0,
    output      wire                                CDOVALID_X0_Y0_D0,
    input       wire                                CDOREADY_X0_Y0_D0,

    //router1
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X0_Y1_D0,
    input       wire                                CDIVALID_X0_Y1_D0,
    output      wire                                CDIREADY_X0_Y1_D0,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X0_Y1_D0,
    output      wire                                CDOVALID_X0_Y1_D0,
    input       wire                                CDOREADY_X0_Y1_D0,

    //router2
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X0_Y2_D0,
    input       wire                                CDIVALID_X0_Y2_D0,
    output      wire                                CDIREADY_X0_Y2_D0,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X0_Y2_D0,
    output      wire                                CDOVALID_X0_Y2_D0,
    input       wire                                CDOREADY_X0_Y2_D0,

    //router3
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X0_Y3_D0,
    input       wire                                CDIVALID_X0_Y3_D0,
    output      wire                                CDIREADY_X0_Y3_D0,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X0_Y3_D0,
    output      wire                                CDOVALID_X0_Y3_D0,
    input       wire                                CDOREADY_X0_Y3_D0,

    //router4
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X0_Y4_D0,
    input       wire                                CDIVALID_X0_Y4_D0,
    output      wire                                CDIREADY_X0_Y4_D0,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X0_Y4_D0,
    output      wire                                CDOVALID_X0_Y4_D0,
    input       wire                                CDOREADY_X0_Y4_D0,

    //router5
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X1_Y0_D0,
    input       wire                                CDIVALID_X1_Y0_D0,
    output      wire                                CDIREADY_X1_Y0_D0,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X1_Y0_D0,
    output      wire                                CDOVALID_X1_Y0_D0,
    input       wire                                CDOREADY_X1_Y0_D0,

    //router6
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X1_Y1_D0,
    input       wire                                CDIVALID_X1_Y1_D0,
    output      wire                                CDIREADY_X1_Y1_D0,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X1_Y1_D0,
    output      wire                                CDOVALID_X1_Y1_D0,
    input       wire                                CDOREADY_X1_Y1_D0,

    //router7
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X1_Y2_D0,
    input       wire                                CDIVALID_X1_Y2_D0,
    output      wire                                CDIREADY_X1_Y2_D0,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X1_Y2_D0,
    output      wire                                CDOVALID_X1_Y2_D0,
    input       wire                                CDOREADY_X1_Y2_D0,

    //router8
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X1_Y3_D0,
    input       wire                                CDIVALID_X1_Y3_D0,
    output      wire                                CDIREADY_X1_Y3_D0,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X1_Y3_D0,
    output      wire                                CDOVALID_X1_Y3_D0,
    input       wire                                CDOREADY_X1_Y3_D0,

    //router9
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X1_Y4_D0,
    input       wire                                CDIVALID_X1_Y4_D0,
    output      wire                                CDIREADY_X1_Y4_D0,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X1_Y4_D0,
    output      wire                                CDOVALID_X1_Y4_D0,
    input       wire                                CDOREADY_X1_Y4_D0,

    // //router10
    // input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X2_Y0,
    // input       wire                                CDIVALID_X2_Y0,
    // output      wire                                CDIREADY_X2_Y0,

    // output      wire        [`DATA_WIDTH-1:0]       CDODATA_X2_Y0,
    // output      wire                                CDOVALID_X2_Y0,
    // input       wire                                CDOREADY_X2_Y0,

    //router11
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X2_Y1_D0,
    input       wire                                CDIVALID_X2_Y1_D0,
    output      wire                                CDIREADY_X2_Y1_D0,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X2_Y1_D0,
    output      wire                                CDOVALID_X2_Y1_D0,
    input       wire                                CDOREADY_X2_Y1_D0,

    //router12
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X2_Y2_D0,
    input       wire                                CDIVALID_X2_Y2_D0,
    output      wire                                CDIREADY_X2_Y2_D0,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X2_Y2_D0,
    output      wire                                CDOVALID_X2_Y2_D0,
    input       wire                                CDOREADY_X2_Y2_D0,

    //router13
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X2_Y3_D0,
    input       wire                                CDIVALID_X2_Y3_D0,
    output      wire                                CDIREADY_X2_Y3_D0,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X2_Y3_D0,
    output      wire                                CDOVALID_X2_Y3_D0,
    input       wire                                CDOREADY_X2_Y3_D0,

    // //router14
    // input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X2_Y4,
    // input       wire                                CDIVALID_X2_Y4,
    // output      wire                                CDIREADY_X2_Y4,

    // output      wire        [`DATA_WIDTH-1:0]       CDODATA_X2_Y4,
    // output      wire                                CDOVALID_X2_Y4,
    // input       wire                                CDOREADY_X2_Y4,

    //router15
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X3_Y0_D0,
    input       wire                                CDIVALID_X3_Y0_D0,
    output      wire                                CDIREADY_X3_Y0_D0,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X3_Y0_D0,
    output      wire                                CDOVALID_X3_Y0_D0,
    input       wire                                CDOREADY_X3_Y0_D0,

    //router16
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X3_Y1_D0,
    input       wire                                CDIVALID_X3_Y1_D0,
    output      wire                                CDIREADY_X3_Y1_D0,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X3_Y1_D0,
    output      wire                                CDOVALID_X3_Y1_D0,
    input       wire                                CDOREADY_X3_Y1_D0,

    //router17
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X3_Y2_D0,
    input       wire                                CDIVALID_X3_Y2_D0,
    output      wire                                CDIREADY_X3_Y2_D0,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X3_Y2_D0,
    output      wire                                CDOVALID_X3_Y2_D0,
    input       wire                                CDOREADY_X3_Y2_D0,

    //router18
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X3_Y3_D0,
    input       wire                                CDIVALID_X3_Y3_D0,
    output      wire                                CDIREADY_X3_Y3_D0,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X3_Y3_D0,
    output      wire                                CDOVALID_X3_Y3_D0,
    input       wire                                CDOREADY_X3_Y3_D0,

    //router19
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X3_Y4_D0,
    input       wire                                CDIVALID_X3_Y4_D0,
    output      wire                                CDIREADY_X3_Y4_D0,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X3_Y4_D0,
    output      wire                                CDOVALID_X3_Y4_D0,
    input       wire                                CDOREADY_X3_Y4_D0,

    //router20
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X4_Y0_D0,
    input       wire                                CDIVALID_X4_Y0_D0,
    output      wire                                CDIREADY_X4_Y0_D0,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X4_Y0_D0,
    output      wire                                CDOVALID_X4_Y0_D0,
    input       wire                                CDOREADY_X4_Y0_D0,

    //router21
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X4_Y1_D0,
    input       wire                                CDIVALID_X4_Y1_D0,
    output      wire                                CDIREADY_X4_Y1_D0,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X4_Y1_D0,
    output      wire                                CDOVALID_X4_Y1_D0,
    input       wire                                CDOREADY_X4_Y1_D0,

    //router22
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X4_Y2_D0,
    input       wire                                CDIVALID_X4_Y2_D0,
    output      wire                                CDIREADY_X4_Y2_D0,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X4_Y2_D0,
    output      wire                                CDOVALID_X4_Y2_D0,
    input       wire                                CDOREADY_X4_Y2_D0,

    //router23
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X4_Y3_D0,
    input       wire                                CDIVALID_X4_Y3_D0,
    output      wire                                CDIREADY_X4_Y3_D0,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X4_Y3_D0,
    output      wire                                CDOVALID_X4_Y3_D0,
    input       wire                                CDOREADY_X4_Y3_D0,

    //router24
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X4_Y4_D0,
    input       wire                                CDIVALID_X4_Y4_D0,
    output      wire                                CDIREADY_X4_Y4_D0,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X4_Y4_D0,
    output      wire                                CDOVALID_X4_Y4_D0,
    input       wire                                CDOREADY_X4_Y4_D0,

    //==============================================================//
    //                                                              /
    //                           NoD1                               /
    //                                                              /
    //==============================================================//
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X0_Y0_D1,
    input       wire                                CDIVALID_X0_Y0_D1,
    output      wire                                CDIREADY_X0_Y0_D1,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X0_Y0_D1,
    output      wire                                CDOVALID_X0_Y0_D1,
    input       wire                                CDOREADY_X0_Y0_D1,

    //router1
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X0_Y1_D1,
    input       wire                                CDIVALID_X0_Y1_D1,
    output      wire                                CDIREADY_X0_Y1_D1,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X0_Y1_D1,
    output      wire                                CDOVALID_X0_Y1_D1,
    input       wire                                CDOREADY_X0_Y1_D1,

    //router2
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X0_Y2_D1,
    input       wire                                CDIVALID_X0_Y2_D1,
    output      wire                                CDIREADY_X0_Y2_D1,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X0_Y2_D1,
    output      wire                                CDOVALID_X0_Y2_D1,
    input       wire                                CDOREADY_X0_Y2_D1,

    //router3
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X0_Y3_D1,
    input       wire                                CDIVALID_X0_Y3_D1,
    output      wire                                CDIREADY_X0_Y3_D1,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X0_Y3_D1,
    output      wire                                CDOVALID_X0_Y3_D1,
    input       wire                                CDOREADY_X0_Y3_D1,

    //router4
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X0_Y4_D1,
    input       wire                                CDIVALID_X0_Y4_D1,
    output      wire                                CDIREADY_X0_Y4_D1,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X0_Y4_D1,
    output      wire                                CDOVALID_X0_Y4_D1,
    input       wire                                CDOREADY_X0_Y4_D1,

    //router5
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X1_Y0_D1,
    input       wire                                CDIVALID_X1_Y0_D1,
    output      wire                                CDIREADY_X1_Y0_D1,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X1_Y0_D1,
    output      wire                                CDOVALID_X1_Y0_D1,
    input       wire                                CDOREADY_X1_Y0_D1,

    //router6
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X1_Y1_D1,
    input       wire                                CDIVALID_X1_Y1_D1,
    output      wire                                CDIREADY_X1_Y1_D1,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X1_Y1_D1,
    output      wire                                CDOVALID_X1_Y1_D1,
    input       wire                                CDOREADY_X1_Y1_D1,

    //router7
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X1_Y2_D1,
    input       wire                                CDIVALID_X1_Y2_D1,
    output      wire                                CDIREADY_X1_Y2_D1,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X1_Y2_D1,
    output      wire                                CDOVALID_X1_Y2_D1,
    input       wire                                CDOREADY_X1_Y2_D1,

    //router8
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X1_Y3_D1,
    input       wire                                CDIVALID_X1_Y3_D1,
    output      wire                                CDIREADY_X1_Y3_D1,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X1_Y3_D1,
    output      wire                                CDOVALID_X1_Y3_D1,
    input       wire                                CDOREADY_X1_Y3_D1,

    //router9
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X1_Y4_D1,
    input       wire                                CDIVALID_X1_Y4_D1,
    output      wire                                CDIREADY_X1_Y4_D1,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X1_Y4_D1,
    output      wire                                CDOVALID_X1_Y4_D1,
    input       wire                                CDOREADY_X1_Y4_D1,

    // //router10
    // input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X2_Y0,
    // input       wire                                CDIVALID_X2_Y0,
    // output      wire                                CDIREADY_X2_Y0,

    // output      wire        [`DATA_WIDTH-1:0]       CDODATA_X2_Y0,
    // output      wire                                CDOVALID_X2_Y0,
    // input       wire                                CDOREADY_X2_Y0,

    //router11
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X2_Y1_D1,
    input       wire                                CDIVALID_X2_Y1_D1,
    output      wire                                CDIREADY_X2_Y1_D1,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X2_Y1_D1,
    output      wire                                CDOVALID_X2_Y1_D1,
    input       wire                                CDOREADY_X2_Y1_D1,

    //router12
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X2_Y2_D1,
    input       wire                                CDIVALID_X2_Y2_D1,
    output      wire                                CDIREADY_X2_Y2_D1,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X2_Y2_D1,
    output      wire                                CDOVALID_X2_Y2_D1,
    input       wire                                CDOREADY_X2_Y2_D1,

    //router13
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X2_Y3_D1,
    input       wire                                CDIVALID_X2_Y3_D1,
    output      wire                                CDIREADY_X2_Y3_D1,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X2_Y3_D1,
    output      wire                                CDOVALID_X2_Y3_D1,
    input       wire                                CDOREADY_X2_Y3_D1,

    // //router14
    // input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X2_Y4,
    // input       wire                                CDIVALID_X2_Y4,
    // output      wire                                CDIREADY_X2_Y4,

    // output      wire        [`DATA_WIDTH-1:0]       CDODATA_X2_Y4,
    // output      wire                                CDOVALID_X2_Y4,
    // input       wire                                CDOREADY_X2_Y4,

    //router15
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X3_Y0_D1,
    input       wire                                CDIVALID_X3_Y0_D1,
    output      wire                                CDIREADY_X3_Y0_D1,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X3_Y0_D1,
    output      wire                                CDOVALID_X3_Y0_D1,
    input       wire                                CDOREADY_X3_Y0_D1,

    //router16
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X3_Y1_D1,
    input       wire                                CDIVALID_X3_Y1_D1,
    output      wire                                CDIREADY_X3_Y1_D1,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X3_Y1_D1,
    output      wire                                CDOVALID_X3_Y1_D1,
    input       wire                                CDOREADY_X3_Y1_D1,

    //router17
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X3_Y2_D1,
    input       wire                                CDIVALID_X3_Y2_D1,
    output      wire                                CDIREADY_X3_Y2_D1,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X3_Y2_D1,
    output      wire                                CDOVALID_X3_Y2_D1,
    input       wire                                CDOREADY_X3_Y2_D1,

    //router18
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X3_Y3_D1,
    input       wire                                CDIVALID_X3_Y3_D1,
    output      wire                                CDIREADY_X3_Y3_D1,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X3_Y3_D1,
    output      wire                                CDOVALID_X3_Y3_D1,
    input       wire                                CDOREADY_X3_Y3_D1,

    //router19
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X3_Y4_D1,
    input       wire                                CDIVALID_X3_Y4_D1,
    output      wire                                CDIREADY_X3_Y4_D1,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X3_Y4_D1,
    output      wire                                CDOVALID_X3_Y4_D1,
    input       wire                                CDOREADY_X3_Y4_D1,

    //router20
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X4_Y0_D1,
    input       wire                                CDIVALID_X4_Y0_D1,
    output      wire                                CDIREADY_X4_Y0_D1,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X4_Y0_D1,
    output      wire                                CDOVALID_X4_Y0_D1,
    input       wire                                CDOREADY_X4_Y0_D1,

    //router21
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X4_Y1_D1,
    input       wire                                CDIVALID_X4_Y1_D1,
    output      wire                                CDIREADY_X4_Y1_D1,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X4_Y1_D1,
    output      wire                                CDOVALID_X4_Y1_D1,
    input       wire                                CDOREADY_X4_Y1_D1,

    //router22
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X4_Y2_D1,
    input       wire                                CDIVALID_X4_Y2_D1,
    output      wire                                CDIREADY_X4_Y2_D1,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X4_Y2_D1,
    output      wire                                CDOVALID_X4_Y2_D1,
    input       wire                                CDOREADY_X4_Y2_D1,

    //router23
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X4_Y3_D1,
    input       wire                                CDIVALID_X4_Y3_D1,
    output      wire                                CDIREADY_X4_Y3_D1,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X4_Y3_D1,
    output      wire                                CDOVALID_X4_Y3_D1,
    input       wire                                CDOREADY_X4_Y3_D1,

    //router24
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X4_Y4_D1,
    input       wire                                CDIVALID_X4_Y4_D1,
    output      wire                                CDIREADY_X4_Y4_D1,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X4_Y4_D1,
    output      wire                                CDOVALID_X4_Y4_D1,
    input       wire                                CDOREADY_X4_Y4_D1,


    //==============================================================//
    //                                                              /
    //                           NoD2                               /
    //                                                              /
    //==============================================================//
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X0_Y0_D2,
    input       wire                                CDIVALID_X0_Y0_D2,
    output      wire                                CDIREADY_X0_Y0_D2,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X0_Y0_D2,
    output      wire                                CDOVALID_X0_Y0_D2,
    input       wire                                CDOREADY_X0_Y0_D2,

    //router1
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X0_Y1_D2,
    input       wire                                CDIVALID_X0_Y1_D2,
    output      wire                                CDIREADY_X0_Y1_D2,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X0_Y1_D2,
    output      wire                                CDOVALID_X0_Y1_D2,
    input       wire                                CDOREADY_X0_Y1_D2,

    //router2
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X0_Y2_D2,
    input       wire                                CDIVALID_X0_Y2_D2,
    output      wire                                CDIREADY_X0_Y2_D2,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X0_Y2_D2,
    output      wire                                CDOVALID_X0_Y2_D2,
    input       wire                                CDOREADY_X0_Y2_D2,

    //router3
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X0_Y3_D2,
    input       wire                                CDIVALID_X0_Y3_D2,
    output      wire                                CDIREADY_X0_Y3_D2,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X0_Y3_D2,
    output      wire                                CDOVALID_X0_Y3_D2,
    input       wire                                CDOREADY_X0_Y3_D2,

    //router4
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X0_Y4_D2,
    input       wire                                CDIVALID_X0_Y4_D2,
    output      wire                                CDIREADY_X0_Y4_D2,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X0_Y4_D2,
    output      wire                                CDOVALID_X0_Y4_D2,
    input       wire                                CDOREADY_X0_Y4_D2,

    //router5
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X1_Y0_D2,
    input       wire                                CDIVALID_X1_Y0_D2,
    output      wire                                CDIREADY_X1_Y0_D2,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X1_Y0_D2,
    output      wire                                CDOVALID_X1_Y0_D2,
    input       wire                                CDOREADY_X1_Y0_D2,

    //router6
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X1_Y1_D2,
    input       wire                                CDIVALID_X1_Y1_D2,
    output      wire                                CDIREADY_X1_Y1_D2,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X1_Y1_D2,
    output      wire                                CDOVALID_X1_Y1_D2,
    input       wire                                CDOREADY_X1_Y1_D2,

    //router7
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X1_Y2_D2,
    input       wire                                CDIVALID_X1_Y2_D2,
    output      wire                                CDIREADY_X1_Y2_D2,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X1_Y2_D2,
    output      wire                                CDOVALID_X1_Y2_D2,
    input       wire                                CDOREADY_X1_Y2_D2,

    //router8
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X1_Y3_D2,
    input       wire                                CDIVALID_X1_Y3_D2,
    output      wire                                CDIREADY_X1_Y3_D2,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X1_Y3_D2,
    output      wire                                CDOVALID_X1_Y3_D2,
    input       wire                                CDOREADY_X1_Y3_D2,

    //router9
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X1_Y4_D2,
    input       wire                                CDIVALID_X1_Y4_D2,
    output      wire                                CDIREADY_X1_Y4_D2,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X1_Y4_D2,
    output      wire                                CDOVALID_X1_Y4_D2,
    input       wire                                CDOREADY_X1_Y4_D2,

    // //router10
    // input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X2_Y0,
    // input       wire                                CDIVALID_X2_Y0,
    // output      wire                                CDIREADY_X2_Y0,

    // output      wire        [`DATA_WIDTH-1:0]       CDODATA_X2_Y0,
    // output      wire                                CDOVALID_X2_Y0,
    // input       wire                                CDOREADY_X2_Y0,

    //router11
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X2_Y1_D2,
    input       wire                                CDIVALID_X2_Y1_D2,
    output      wire                                CDIREADY_X2_Y1_D2,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X2_Y1_D2,
    output      wire                                CDOVALID_X2_Y1_D2,
    input       wire                                CDOREADY_X2_Y1_D2,

    //router12
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X2_Y2_D2,
    input       wire                                CDIVALID_X2_Y2_D2,
    output      wire                                CDIREADY_X2_Y2_D2,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X2_Y2_D2,
    output      wire                                CDOVALID_X2_Y2_D2,
    input       wire                                CDOREADY_X2_Y2_D2,

    //router13
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X2_Y3_D2,
    input       wire                                CDIVALID_X2_Y3_D2,
    output      wire                                CDIREADY_X2_Y3_D2,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X2_Y3_D2,
    output      wire                                CDOVALID_X2_Y3_D2,
    input       wire                                CDOREADY_X2_Y3_D2,

    // //router14
    // input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X2_Y4,
    // input       wire                                CDIVALID_X2_Y4,
    // output      wire                                CDIREADY_X2_Y4,

    // output      wire        [`DATA_WIDTH-1:0]       CDODATA_X2_Y4,
    // output      wire                                CDOVALID_X2_Y4,
    // input       wire                                CDOREADY_X2_Y4,

    //router15
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X3_Y0_D2,
    input       wire                                CDIVALID_X3_Y0_D2,
    output      wire                                CDIREADY_X3_Y0_D2,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X3_Y0_D2,
    output      wire                                CDOVALID_X3_Y0_D2,
    input       wire                                CDOREADY_X3_Y0_D2,

    //router16
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X3_Y1_D2,
    input       wire                                CDIVALID_X3_Y1_D2,
    output      wire                                CDIREADY_X3_Y1_D2,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X3_Y1_D2,
    output      wire                                CDOVALID_X3_Y1_D2,
    input       wire                                CDOREADY_X3_Y1_D2,

    //router17
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X3_Y2_D2,
    input       wire                                CDIVALID_X3_Y2_D2,
    output      wire                                CDIREADY_X3_Y2_D2,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X3_Y2_D2,
    output      wire                                CDOVALID_X3_Y2_D2,
    input       wire                                CDOREADY_X3_Y2_D2,

    //router18
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X3_Y3_D2,
    input       wire                                CDIVALID_X3_Y3_D2,
    output      wire                                CDIREADY_X3_Y3_D2,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X3_Y3_D2,
    output      wire                                CDOVALID_X3_Y3_D2,
    input       wire                                CDOREADY_X3_Y3_D2,

    //router19
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X3_Y4_D2,
    input       wire                                CDIVALID_X3_Y4_D2,
    output      wire                                CDIREADY_X3_Y4_D2,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X3_Y4_D2,
    output      wire                                CDOVALID_X3_Y4_D2,
    input       wire                                CDOREADY_X3_Y4_D2,

    //router20
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X4_Y0_D2,
    input       wire                                CDIVALID_X4_Y0_D2,
    output      wire                                CDIREADY_X4_Y0_D2,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X4_Y0_D2,
    output      wire                                CDOVALID_X4_Y0_D2,
    input       wire                                CDOREADY_X4_Y0_D2,

    //router21
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X4_Y1_D2,
    input       wire                                CDIVALID_X4_Y1_D2,
    output      wire                                CDIREADY_X4_Y1_D2,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X4_Y1_D2,
    output      wire                                CDOVALID_X4_Y1_D2,
    input       wire                                CDOREADY_X4_Y1_D2,

    //router22
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X4_Y2_D2,
    input       wire                                CDIVALID_X4_Y2_D2,
    output      wire                                CDIREADY_X4_Y2_D2,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X4_Y2_D2,
    output      wire                                CDOVALID_X4_Y2_D2,
    input       wire                                CDOREADY_X4_Y2_D2,

    //router23
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X4_Y3_D2,
    input       wire                                CDIVALID_X4_Y3_D2,
    output      wire                                CDIREADY_X4_Y3_D2,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X4_Y3_D2,
    output      wire                                CDOVALID_X4_Y3_D2,
    input       wire                                CDOREADY_X4_Y3_D2,

    //router24
    input       wire        [`DATA_WIDTH-1:0]       CDIDATA_X4_Y4_D2,
    input       wire                                CDIVALID_X4_Y4_D2,
    output      wire                                CDIREADY_X4_Y4_D2,

    output      wire        [`DATA_WIDTH-1:0]       CDODATA_X4_Y4_D2,
    output      wire                                CDOVALID_X4_Y4_D2,
    input       wire                                CDOREADY_X4_Y4_D2
);

wire [`DATA_WIDTH/2-1:0] d0_2_d1_data,d1_2_d0_data,d1_2_d2_data,d2_2_d1_data;
wire d0_2_d1_valid,d1_2_d0_valid,d1_2_d2_valid,d2_2_d1_valid;
wire d0_2_d1_ready,d1_2_d0_ready,d1_2_d2_ready,d2_2_d1_ready;

ExtenNoD #(
    .NODID                        (0)
)NoD0(
    .CDCLK                        (CDCLK),
    .CPCLK                        (CPCLK),
    .CDRESETn                     (CDRESETn),
    .CDIDATA_X0_Y0                (CDIDATA_X0_Y0_D0), 
    .CDIVALID_X0_Y0               (CDIVALID_X0_Y0_D0),
    .CDIREADY_X0_Y0               (CDIREADY_X0_Y0_D0),
    .CDODATA_X0_Y0                (CDODATA_X0_Y0_D0), 
    .CDOVALID_X0_Y0               (CDOVALID_X0_Y0_D0),
    .CDOREADY_X0_Y0               (CDOREADY_X0_Y0_D0),
    .CDIDATA_X0_Y1                (CDIDATA_X0_Y1_D0), 
    .CDIVALID_X0_Y1               (CDIVALID_X0_Y1_D0),
    .CDIREADY_X0_Y1               (CDIREADY_X0_Y1_D0),
    .CDODATA_X0_Y1                (CDODATA_X0_Y1_D0), 
    .CDOVALID_X0_Y1               (CDOVALID_X0_Y1_D0),
    .CDOREADY_X0_Y1               (CDOREADY_X0_Y1_D0),
    .CDIDATA_X0_Y2                (CDIDATA_X0_Y2_D0), 
    .CDIVALID_X0_Y2               (CDIVALID_X0_Y2_D0),
    .CDIREADY_X0_Y2               (CDIREADY_X0_Y2_D0),
    .CDODATA_X0_Y2                (CDODATA_X0_Y2_D0), 
    .CDOVALID_X0_Y2               (CDOVALID_X0_Y2_D0),
    .CDOREADY_X0_Y2               (CDOREADY_X0_Y2_D0),
    .CDIDATA_X0_Y3                (CDIDATA_X0_Y3_D0), 
    .CDIVALID_X0_Y3               (CDIVALID_X0_Y3_D0),
    .CDIREADY_X0_Y3               (CDIREADY_X0_Y3_D0),
    .CDODATA_X0_Y3                (CDODATA_X0_Y3_D0),
    .CDOVALID_X0_Y3               (CDOVALID_X0_Y3_D0),
    .CDOREADY_X0_Y3               (CDOREADY_X0_Y3_D0),
    .CDIDATA_X0_Y4                (CDIDATA_X0_Y4_D0),
    .CDIVALID_X0_Y4               (CDIVALID_X0_Y4_D0),
    .CDIREADY_X0_Y4               (CDIREADY_X0_Y4_D0),
    .CDODATA_X0_Y4                (CDODATA_X0_Y4_D0),
    .CDOVALID_X0_Y4               (CDOVALID_X0_Y4_D0),
    .CDOREADY_X0_Y4               (CDOREADY_X0_Y4_D0),
    .CDIDATA_X1_Y0                (CDIDATA_X1_Y0_D0),
    .CDIVALID_X1_Y0               (CDIVALID_X1_Y0_D0),
    .CDIREADY_X1_Y0               (CDIREADY_X1_Y0_D0),
    .CDODATA_X1_Y0                (CDODATA_X1_Y0_D0),
    .CDOVALID_X1_Y0               (CDOVALID_X1_Y0_D0),
    .CDOREADY_X1_Y0               (CDOREADY_X1_Y0_D0),
    .CDIDATA_X1_Y1                (CDIDATA_X1_Y1_D0),
    .CDIVALID_X1_Y1               (CDIVALID_X1_Y1_D0),
    .CDIREADY_X1_Y1               (CDIREADY_X1_Y1_D0),
    .CDODATA_X1_Y1                (CDODATA_X1_Y1_D0),
    .CDOVALID_X1_Y1               (CDOVALID_X1_Y1_D0),
    .CDOREADY_X1_Y1               (CDOREADY_X1_Y1_D0),
    .CDIDATA_X1_Y2                (CDIDATA_X1_Y2_D0),
    .CDIVALID_X1_Y2               (CDIVALID_X1_Y2_D0),
    .CDIREADY_X1_Y2               (CDIREADY_X1_Y2_D0),
    .CDODATA_X1_Y2                (CDODATA_X1_Y2_D0),
    .CDOVALID_X1_Y2               (CDOVALID_X1_Y2_D0),
    .CDOREADY_X1_Y2               (CDOREADY_X1_Y2_D0),
    .CDIDATA_X1_Y3                (CDIDATA_X1_Y3_D0),
    .CDIVALID_X1_Y3               (CDIVALID_X1_Y3_D0),
    .CDIREADY_X1_Y3               (CDIREADY_X1_Y3_D0),
    .CDODATA_X1_Y3                (CDODATA_X1_Y3_D0),
    .CDOVALID_X1_Y3               (CDOVALID_X1_Y3_D0),
    .CDOREADY_X1_Y3               (CDOREADY_X1_Y3_D0),
    .CDIDATA_X1_Y4                (CDIDATA_X1_Y4_D0),
    .CDIVALID_X1_Y4               (CDIVALID_X1_Y4_D0),
    .CDIREADY_X1_Y4               (CDIREADY_X1_Y4_D0),
    .CDODATA_X1_Y4                (CDODATA_X1_Y4_D0),
    .CDOVALID_X1_Y4               (CDOVALID_X1_Y4_D0),
    .CDOREADY_X1_Y4               (CDOREADY_X1_Y4_D0),
    .CDIDATA_X2_Y1                (CDIDATA_X2_Y1_D0),
    .CDIVALID_X2_Y1               (CDIVALID_X2_Y1_D0),
    .CDIREADY_X2_Y1               (CDIREADY_X2_Y1_D0),
    .CDODATA_X2_Y1                (CDODATA_X2_Y1_D0),
    .CDOVALID_X2_Y1               (CDOVALID_X2_Y1_D0),
    .CDOREADY_X2_Y1               (CDOREADY_X2_Y1_D0),
    .CDIDATA_X2_Y2                (CDIDATA_X2_Y2_D0),
    .CDIVALID_X2_Y2               (CDIVALID_X2_Y2_D0),
    .CDIREADY_X2_Y2               (CDIREADY_X2_Y2_D0),
    .CDODATA_X2_Y2                (CDODATA_X2_Y2_D0),
    .CDOVALID_X2_Y2               (CDOVALID_X2_Y2_D0),
    .CDOREADY_X2_Y2               (CDOREADY_X2_Y2_D0),
    .CDIDATA_X2_Y3                (CDIDATA_X2_Y3_D0),
    .CDIVALID_X2_Y3               (CDIVALID_X2_Y3_D0),
    .CDIREADY_X2_Y3               (CDIREADY_X2_Y3_D0),
    .CDODATA_X2_Y3                (CDODATA_X2_Y3_D0),
    .CDOVALID_X2_Y3               (CDOVALID_X2_Y3_D0),
    .CDOREADY_X2_Y3               (CDOREADY_X2_Y3_D0),
    .CDIDATA_X3_Y0                (CDIDATA_X3_Y0_D0),
    .CDIVALID_X3_Y0               (CDIVALID_X3_Y0_D0),
    .CDIREADY_X3_Y0               (CDIREADY_X3_Y0_D0),
    .CDODATA_X3_Y0                (CDODATA_X3_Y0_D0),
    .CDOVALID_X3_Y0               (CDOVALID_X3_Y0_D0),
    .CDOREADY_X3_Y0               (CDOREADY_X3_Y0_D0),
    .CDIDATA_X3_Y1                (CDIDATA_X3_Y1_D0),
    .CDIVALID_X3_Y1               (CDIVALID_X3_Y1_D0),
    .CDIREADY_X3_Y1               (CDIREADY_X3_Y1_D0),
    .CDODATA_X3_Y1                (CDODATA_X3_Y1_D0),
    .CDOVALID_X3_Y1               (CDOVALID_X3_Y1_D0),
    .CDOREADY_X3_Y1               (CDOREADY_X3_Y1_D0),
    .CDIDATA_X3_Y2                (CDIDATA_X3_Y2_D0),
    .CDIVALID_X3_Y2               (CDIVALID_X3_Y2_D0),
    .CDIREADY_X3_Y2               (CDIREADY_X3_Y2_D0),
    .CDODATA_X3_Y2                (CDODATA_X3_Y2_D0),
    .CDOVALID_X3_Y2               (CDOVALID_X3_Y2_D0),
    .CDOREADY_X3_Y2               (CDOREADY_X3_Y2_D0),
    .CDIDATA_X3_Y3                (CDIDATA_X3_Y3_D0),
    .CDIVALID_X3_Y3               (CDIVALID_X3_Y3_D0),
    .CDIREADY_X3_Y3               (CDIREADY_X3_Y3_D0),
    .CDODATA_X3_Y3                (CDODATA_X3_Y3_D0),
    .CDOVALID_X3_Y3               (CDOVALID_X3_Y3_D0),
    .CDOREADY_X3_Y3               (CDOREADY_X3_Y3_D0),
    .CDIDATA_X3_Y4                (CDIDATA_X3_Y4_D0),
    .CDIVALID_X3_Y4               (CDIVALID_X3_Y4_D0),
    .CDIREADY_X3_Y4               (CDIREADY_X3_Y4_D0),
    .CDODATA_X3_Y4                (CDODATA_X3_Y4_D0),
    .CDOVALID_X3_Y4               (CDOVALID_X3_Y4_D0),
    .CDOREADY_X3_Y4               (CDOREADY_X3_Y4_D0),
    .CDIDATA_X4_Y0                (CDIDATA_X4_Y0_D0),
    .CDIVALID_X4_Y0               (CDIVALID_X4_Y0_D0),
    .CDIREADY_X4_Y0               (CDIREADY_X4_Y0_D0),
    .CDODATA_X4_Y0                (CDODATA_X4_Y0_D0),
    .CDOVALID_X4_Y0               (CDOVALID_X4_Y0_D0),
    .CDOREADY_X4_Y0               (CDOREADY_X4_Y0_D0),
    .CDIDATA_X4_Y1                (CDIDATA_X4_Y1_D0),
    .CDIVALID_X4_Y1               (CDIVALID_X4_Y1_D0),
    .CDIREADY_X4_Y1               (CDIREADY_X4_Y1_D0),
    .CDODATA_X4_Y1                (CDODATA_X4_Y1_D0),
    .CDOVALID_X4_Y1               (CDOVALID_X4_Y1_D0),
    .CDOREADY_X4_Y1               (CDOREADY_X4_Y1_D0),
    .CDIDATA_X4_Y2                (CDIDATA_X4_Y2_D0),
    .CDIVALID_X4_Y2               (CDIVALID_X4_Y2_D0),
    .CDIREADY_X4_Y2               (CDIREADY_X4_Y2_D0),
    .CDODATA_X4_Y2                (CDODATA_X4_Y2_D0),
    .CDOVALID_X4_Y2               (CDOVALID_X4_Y2_D0),
    .CDOREADY_X4_Y2               (CDOREADY_X4_Y2_D0),
    .CDIDATA_X4_Y3                (CDIDATA_X4_Y3_D0),
    .CDIVALID_X4_Y3               (CDIVALID_X4_Y3_D0),
    .CDIREADY_X4_Y3               (CDIREADY_X4_Y3_D0),
    .CDODATA_X4_Y3                (CDODATA_X4_Y3_D0),
    .CDOVALID_X4_Y3               (CDOVALID_X4_Y3_D0),
    .CDOREADY_X4_Y3               (CDOREADY_X4_Y3_D0),
    .CDIDATA_X4_Y4                (CDIDATA_X4_Y4_D0),
    .CDIVALID_X4_Y4               (CDIVALID_X4_Y4_D0),
    .CDIREADY_X4_Y4               (CDIREADY_X4_Y4_D0),
    .CDODATA_X4_Y4                (CDODATA_X4_Y4_D0),
    .CDOVALID_X4_Y4               (CDOVALID_X4_Y4_D0),
    .CDOREADY_X4_Y4               (CDOREADY_X4_Y4_D0),
    .CPIDATA_W                    (65'b0),
    .CPIVALID_W                   (1'b0),
    .CPIREADY_W                   (),
    .CPODATA_W                    (),
    .CPOVALID_W                   (),
    .CPOREADY_W                   (1'b0),
    .CPIDATA_E                    (d1_2_d0_data),
    .CPIVALID_E                   (d1_2_d0_valid),
    .CPIREADY_E                   (d1_2_d0_ready),
    .CPODATA_E                    (d0_2_d1_data),
    .CPOVALID_E                   (d0_2_d1_valid),
    .CPOREADY_E                   (d0_2_d1_ready)
);

ExtenNoD #(
    .NODID                        (1)
)NoD1(
    .CDCLK                        (CDCLK),
    .CPCLK                        (CPCLK),
    .CDRESETn                     (CDRESETn),
    .CDIDATA_X0_Y0                (CDIDATA_X0_Y0_D1),
    .CDIVALID_X0_Y0               (CDIVALID_X0_Y0_D1),
    .CDIREADY_X0_Y0               (CDIREADY_X0_Y0_D1),
    .CDODATA_X0_Y0                (CDODATA_X0_Y0_D1),
    .CDOVALID_X0_Y0               (CDOVALID_X0_Y0_D1),
    .CDOREADY_X0_Y0               (CDOREADY_X0_Y0_D1),
    .CDIDATA_X0_Y1                (CDIDATA_X0_Y1_D1),
    .CDIVALID_X0_Y1               (CDIVALID_X0_Y1_D1),
    .CDIREADY_X0_Y1               (CDIREADY_X0_Y1_D1),
    .CDODATA_X0_Y1                (CDODATA_X0_Y1_D1),
    .CDOVALID_X0_Y1               (CDOVALID_X0_Y1_D1),
    .CDOREADY_X0_Y1               (CDOREADY_X0_Y1_D1),
    .CDIDATA_X0_Y2                (CDIDATA_X0_Y2_D1),
    .CDIVALID_X0_Y2               (CDIVALID_X0_Y2_D1),
    .CDIREADY_X0_Y2               (CDIREADY_X0_Y2_D1),
    .CDODATA_X0_Y2                (CDODATA_X0_Y2_D1),
    .CDOVALID_X0_Y2               (CDOVALID_X0_Y2_D1),
    .CDOREADY_X0_Y2               (CDOREADY_X0_Y2_D1),
    .CDIDATA_X0_Y3                (CDIDATA_X0_Y3_D1),
    .CDIVALID_X0_Y3               (CDIVALID_X0_Y3_D1),
    .CDIREADY_X0_Y3               (CDIREADY_X0_Y3_D1),
    .CDODATA_X0_Y3                (CDODATA_X0_Y3_D1),
    .CDOVALID_X0_Y3               (CDOVALID_X0_Y3_D1),
    .CDOREADY_X0_Y3               (CDOREADY_X0_Y3_D1),
    .CDIDATA_X0_Y4                (CDIDATA_X0_Y4_D1),
    .CDIVALID_X0_Y4               (CDIVALID_X0_Y4_D1),
    .CDIREADY_X0_Y4               (CDIREADY_X0_Y4_D1),
    .CDODATA_X0_Y4                (CDODATA_X0_Y4_D1),
    .CDOVALID_X0_Y4               (CDOVALID_X0_Y4_D1),
    .CDOREADY_X0_Y4               (CDOREADY_X0_Y4_D1),
    .CDIDATA_X1_Y0                (CDIDATA_X1_Y0_D1),
    .CDIVALID_X1_Y0               (CDIVALID_X1_Y0_D1),
    .CDIREADY_X1_Y0               (CDIREADY_X1_Y0_D1),
    .CDODATA_X1_Y0                (CDODATA_X1_Y0_D1),
    .CDOVALID_X1_Y0               (CDOVALID_X1_Y0_D1),
    .CDOREADY_X1_Y0               (CDOREADY_X1_Y0_D1),
    .CDIDATA_X1_Y1                (CDIDATA_X1_Y1_D1),
    .CDIVALID_X1_Y1               (CDIVALID_X1_Y1_D1),
    .CDIREADY_X1_Y1               (CDIREADY_X1_Y1_D1),
    .CDODATA_X1_Y1                (CDODATA_X1_Y1_D1),
    .CDOVALID_X1_Y1               (CDOVALID_X1_Y1_D1),
    .CDOREADY_X1_Y1               (CDOREADY_X1_Y1_D1),
    .CDIDATA_X1_Y2                (CDIDATA_X1_Y2_D1),
    .CDIVALID_X1_Y2               (CDIVALID_X1_Y2_D1),
    .CDIREADY_X1_Y2               (CDIREADY_X1_Y2_D1),
    .CDODATA_X1_Y2                (CDODATA_X1_Y2_D1),
    .CDOVALID_X1_Y2               (CDOVALID_X1_Y2_D1),
    .CDOREADY_X1_Y2               (CDOREADY_X1_Y2_D1),
    .CDIDATA_X1_Y3                (CDIDATA_X1_Y3_D1),
    .CDIVALID_X1_Y3               (CDIVALID_X1_Y3_D1),
    .CDIREADY_X1_Y3               (CDIREADY_X1_Y3_D1),
    .CDODATA_X1_Y3                (CDODATA_X1_Y3_D1),
    .CDOVALID_X1_Y3               (CDOVALID_X1_Y3_D1),
    .CDOREADY_X1_Y3               (CDOREADY_X1_Y3_D1),
    .CDIDATA_X1_Y4                (CDIDATA_X1_Y4_D1),
    .CDIVALID_X1_Y4               (CDIVALID_X1_Y4_D1),
    .CDIREADY_X1_Y4               (CDIREADY_X1_Y4_D1),
    .CDODATA_X1_Y4                (CDODATA_X1_Y4_D1),
    .CDOVALID_X1_Y4               (CDOVALID_X1_Y4_D1),
    .CDOREADY_X1_Y4               (CDOREADY_X1_Y4_D1),
    .CDIDATA_X2_Y1                (CDIDATA_X2_Y1_D1),
    .CDIVALID_X2_Y1               (CDIVALID_X2_Y1_D1),
    .CDIREADY_X2_Y1               (CDIREADY_X2_Y1_D1),
    .CDODATA_X2_Y1                (CDODATA_X2_Y1_D1),
    .CDOVALID_X2_Y1               (CDOVALID_X2_Y1_D1),
    .CDOREADY_X2_Y1               (CDOREADY_X2_Y1_D1),
    .CDIDATA_X2_Y2                (CDIDATA_X2_Y2_D1),
    .CDIVALID_X2_Y2               (CDIVALID_X2_Y2_D1),
    .CDIREADY_X2_Y2               (CDIREADY_X2_Y2_D1),
    .CDODATA_X2_Y2                (CDODATA_X2_Y2_D1),
    .CDOVALID_X2_Y2               (CDOVALID_X2_Y2_D1),
    .CDOREADY_X2_Y2               (CDOREADY_X2_Y2_D1),
    .CDIDATA_X2_Y3                (CDIDATA_X2_Y3_D1),
    .CDIVALID_X2_Y3               (CDIVALID_X2_Y3_D1),
    .CDIREADY_X2_Y3               (CDIREADY_X2_Y3_D1),
    .CDODATA_X2_Y3                (CDODATA_X2_Y3_D1),
    .CDOVALID_X2_Y3               (CDOVALID_X2_Y3_D1),
    .CDOREADY_X2_Y3               (CDOREADY_X2_Y3_D1),
    .CDIDATA_X3_Y0                (CDIDATA_X3_Y0_D1),
    .CDIVALID_X3_Y0               (CDIVALID_X3_Y0_D1),
    .CDIREADY_X3_Y0               (CDIREADY_X3_Y0_D1),
    .CDODATA_X3_Y0                (CDODATA_X3_Y0_D1),
    .CDOVALID_X3_Y0               (CDOVALID_X3_Y0_D1),
    .CDOREADY_X3_Y0               (CDOREADY_X3_Y0_D1),
    .CDIDATA_X3_Y1                (CDIDATA_X3_Y1_D1),
    .CDIVALID_X3_Y1               (CDIVALID_X3_Y1_D1),
    .CDIREADY_X3_Y1               (CDIREADY_X3_Y1_D1),
    .CDODATA_X3_Y1                (CDODATA_X3_Y1_D1),
    .CDOVALID_X3_Y1               (CDOVALID_X3_Y1_D1),
    .CDOREADY_X3_Y1               (CDOREADY_X3_Y1_D1),
    .CDIDATA_X3_Y2                (CDIDATA_X3_Y2_D1),
    .CDIVALID_X3_Y2               (CDIVALID_X3_Y2_D1),
    .CDIREADY_X3_Y2               (CDIREADY_X3_Y2_D1),
    .CDODATA_X3_Y2                (CDODATA_X3_Y2_D1),
    .CDOVALID_X3_Y2               (CDOVALID_X3_Y2_D1),
    .CDOREADY_X3_Y2               (CDOREADY_X3_Y2_D1),
    .CDIDATA_X3_Y3                (CDIDATA_X3_Y3_D1),
    .CDIVALID_X3_Y3               (CDIVALID_X3_Y3_D1),
    .CDIREADY_X3_Y3               (CDIREADY_X3_Y3_D1),
    .CDODATA_X3_Y3                (CDODATA_X3_Y3_D1),
    .CDOVALID_X3_Y3               (CDOVALID_X3_Y3_D1),
    .CDOREADY_X3_Y3               (CDOREADY_X3_Y3_D1),
    .CDIDATA_X3_Y4                (CDIDATA_X3_Y4_D1),
    .CDIVALID_X3_Y4               (CDIVALID_X3_Y4_D1),
    .CDIREADY_X3_Y4               (CDIREADY_X3_Y4_D1),
    .CDODATA_X3_Y4                (CDODATA_X3_Y4_D1),
    .CDOVALID_X3_Y4               (CDOVALID_X3_Y4_D1),
    .CDOREADY_X3_Y4               (CDOREADY_X3_Y4_D1),
    .CDIDATA_X4_Y0                (CDIDATA_X4_Y0_D1),
    .CDIVALID_X4_Y0               (CDIVALID_X4_Y0_D1),
    .CDIREADY_X4_Y0               (CDIREADY_X4_Y0_D1),
    .CDODATA_X4_Y0                (CDODATA_X4_Y0_D1),
    .CDOVALID_X4_Y0               (CDOVALID_X4_Y0_D1),
    .CDOREADY_X4_Y0               (CDOREADY_X4_Y0_D1),
    .CDIDATA_X4_Y1                (CDIDATA_X4_Y1_D1),
    .CDIVALID_X4_Y1               (CDIVALID_X4_Y1_D1),
    .CDIREADY_X4_Y1               (CDIREADY_X4_Y1_D1),
    .CDODATA_X4_Y1                (CDODATA_X4_Y1_D1),
    .CDOVALID_X4_Y1               (CDOVALID_X4_Y1_D1),
    .CDOREADY_X4_Y1               (CDOREADY_X4_Y1_D1),
    .CDIDATA_X4_Y2                (CDIDATA_X4_Y2_D1),
    .CDIVALID_X4_Y2               (CDIVALID_X4_Y2_D1),
    .CDIREADY_X4_Y2               (CDIREADY_X4_Y2_D1),
    .CDODATA_X4_Y2                (CDODATA_X4_Y2_D1),
    .CDOVALID_X4_Y2               (CDOVALID_X4_Y2_D1),
    .CDOREADY_X4_Y2               (CDOREADY_X4_Y2_D1),
    .CDIDATA_X4_Y3                (CDIDATA_X4_Y3_D1),
    .CDIVALID_X4_Y3               (CDIVALID_X4_Y3_D1),
    .CDIREADY_X4_Y3               (CDIREADY_X4_Y3_D1),
    .CDODATA_X4_Y3                (CDODATA_X4_Y3_D1),
    .CDOVALID_X4_Y3               (CDOVALID_X4_Y3_D1),
    .CDOREADY_X4_Y3               (CDOREADY_X4_Y3_D1),
    .CDIDATA_X4_Y4                (CDIDATA_X4_Y4_D1),
    .CDIVALID_X4_Y4               (CDIVALID_X4_Y4_D1),
    .CDIREADY_X4_Y4               (CDIREADY_X4_Y4_D1),
    .CDODATA_X4_Y4                (CDODATA_X4_Y4_D1),
    .CDOVALID_X4_Y4               (CDOVALID_X4_Y4_D1),
    .CDOREADY_X4_Y4               (CDOREADY_X4_Y4_D1),
    .CPIDATA_W                    (d0_2_d1_data),
    .CPIVALID_W                   (d0_2_d1_valid),
    .CPIREADY_W                   (d0_2_d1_ready),
    .CPODATA_W                    (d1_2_d0_data),
    .CPOVALID_W                   (d1_2_d0_valid),
    .CPOREADY_W                   (d1_2_d0_ready),
    .CPIDATA_E                    (d2_2_d1_data),
    .CPIVALID_E                   (d2_2_d1_valid),
    .CPIREADY_E                   (d2_2_d1_ready),
    .CPODATA_E                    (d1_2_d2_data),
    .CPOVALID_E                   (d1_2_d2_valid),
    .CPOREADY_E                   (d1_2_d2_ready)
);

ExtenNoD #(
    .NODID                        (2)
)NoD2(
    .CDCLK                        (CDCLK),
    .CPCLK                        (CPCLK),
    .CDRESETn                     (CDRESETn),
    .CDIDATA_X0_Y0                (CDIDATA_X0_Y0_D2),
    .CDIVALID_X0_Y0               (CDIVALID_X0_Y0_D2),
    .CDIREADY_X0_Y0               (CDIREADY_X0_Y0_D2),
    .CDODATA_X0_Y0                (CDODATA_X0_Y0_D2),
    .CDOVALID_X0_Y0               (CDOVALID_X0_Y0_D2),
    .CDOREADY_X0_Y0               (CDOREADY_X0_Y0_D2),
    .CDIDATA_X0_Y1                (CDIDATA_X0_Y1_D2),
    .CDIVALID_X0_Y1               (CDIVALID_X0_Y1_D2),
    .CDIREADY_X0_Y1               (CDIREADY_X0_Y1_D2),
    .CDODATA_X0_Y1                (CDODATA_X0_Y1_D2),
    .CDOVALID_X0_Y1               (CDOVALID_X0_Y1_D2),
    .CDOREADY_X0_Y1               (CDOREADY_X0_Y1_D2),
    .CDIDATA_X0_Y2                (CDIDATA_X0_Y2_D2),
    .CDIVALID_X0_Y2               (CDIVALID_X0_Y2_D2),
    .CDIREADY_X0_Y2               (CDIREADY_X0_Y2_D2),
    .CDODATA_X0_Y2                (CDODATA_X0_Y2_D2),
    .CDOVALID_X0_Y2               (CDOVALID_X0_Y2_D2),
    .CDOREADY_X0_Y2               (CDOREADY_X0_Y2_D2),
    .CDIDATA_X0_Y3                (CDIDATA_X0_Y3_D2),
    .CDIVALID_X0_Y3               (CDIVALID_X0_Y3_D2),
    .CDIREADY_X0_Y3               (CDIREADY_X0_Y3_D2),
    .CDODATA_X0_Y3                (CDODATA_X0_Y3_D2),
    .CDOVALID_X0_Y3               (CDOVALID_X0_Y3_D2),
    .CDOREADY_X0_Y3               (CDOREADY_X0_Y3_D2),
    .CDIDATA_X0_Y4                (CDIDATA_X0_Y4_D2),
    .CDIVALID_X0_Y4               (CDIVALID_X0_Y4_D2),
    .CDIREADY_X0_Y4               (CDIREADY_X0_Y4_D2),
    .CDODATA_X0_Y4                (CDODATA_X0_Y4_D2),
    .CDOVALID_X0_Y4               (CDOVALID_X0_Y4_D2),
    .CDOREADY_X0_Y4               (CDOREADY_X0_Y4_D2),
    .CDIDATA_X1_Y0                (CDIDATA_X1_Y0_D2),
    .CDIVALID_X1_Y0               (CDIVALID_X1_Y0_D2),
    .CDIREADY_X1_Y0               (CDIREADY_X1_Y0_D2),
    .CDODATA_X1_Y0                (CDODATA_X1_Y0_D2),
    .CDOVALID_X1_Y0               (CDOVALID_X1_Y0_D2),
    .CDOREADY_X1_Y0               (CDOREADY_X1_Y0_D2),
    .CDIDATA_X1_Y1                (CDIDATA_X1_Y1_D2),
    .CDIVALID_X1_Y1               (CDIVALID_X1_Y1_D2),
    .CDIREADY_X1_Y1               (CDIREADY_X1_Y1_D2),
    .CDODATA_X1_Y1                (CDODATA_X1_Y1_D2),
    .CDOVALID_X1_Y1               (CDOVALID_X1_Y1_D2),
    .CDOREADY_X1_Y1               (CDOREADY_X1_Y1_D2),
    .CDIDATA_X1_Y2                (CDIDATA_X1_Y2_D2),
    .CDIVALID_X1_Y2               (CDIVALID_X1_Y2_D2),
    .CDIREADY_X1_Y2               (CDIREADY_X1_Y2_D2),
    .CDODATA_X1_Y2                (CDODATA_X1_Y2_D2),
    .CDOVALID_X1_Y2               (CDOVALID_X1_Y2_D2),
    .CDOREADY_X1_Y2               (CDOREADY_X1_Y2_D2),
    .CDIDATA_X1_Y3                (CDIDATA_X1_Y3_D2),
    .CDIVALID_X1_Y3               (CDIVALID_X1_Y3_D2),
    .CDIREADY_X1_Y3               (CDIREADY_X1_Y3_D2),
    .CDODATA_X1_Y3                (CDODATA_X1_Y3_D2),
    .CDOVALID_X1_Y3               (CDOVALID_X1_Y3_D2),
    .CDOREADY_X1_Y3               (CDOREADY_X1_Y3_D2),
    .CDIDATA_X1_Y4                (CDIDATA_X1_Y4_D2),
    .CDIVALID_X1_Y4               (CDIVALID_X1_Y4_D2),
    .CDIREADY_X1_Y4               (CDIREADY_X1_Y4_D2),
    .CDODATA_X1_Y4                (CDODATA_X1_Y4_D2),
    .CDOVALID_X1_Y4               (CDOVALID_X1_Y4_D2),
    .CDOREADY_X1_Y4               (CDOREADY_X1_Y4_D2),
    .CDIDATA_X2_Y1                (CDIDATA_X2_Y1_D2),
    .CDIVALID_X2_Y1               (CDIVALID_X2_Y1_D2),
    .CDIREADY_X2_Y1               (CDIREADY_X2_Y1_D2),
    .CDODATA_X2_Y1                (CDODATA_X2_Y1_D2),
    .CDOVALID_X2_Y1               (CDOVALID_X2_Y1_D2),
    .CDOREADY_X2_Y1               (CDOREADY_X2_Y1_D2),
    .CDIDATA_X2_Y2                (CDIDATA_X2_Y2_D2),
    .CDIVALID_X2_Y2               (CDIVALID_X2_Y2_D2),
    .CDIREADY_X2_Y2               (CDIREADY_X2_Y2_D2),
    .CDODATA_X2_Y2                (CDODATA_X2_Y2_D2),
    .CDOVALID_X2_Y2               (CDOVALID_X2_Y2_D2),
    .CDOREADY_X2_Y2               (CDOREADY_X2_Y2_D2),
    .CDIDATA_X2_Y3                (CDIDATA_X2_Y3_D2),
    .CDIVALID_X2_Y3               (CDIVALID_X2_Y3_D2),
    .CDIREADY_X2_Y3               (CDIREADY_X2_Y3_D2),
    .CDODATA_X2_Y3                (CDODATA_X2_Y3_D2),
    .CDOVALID_X2_Y3               (CDOVALID_X2_Y3_D2),
    .CDOREADY_X2_Y3               (CDOREADY_X2_Y3_D2),
    .CDIDATA_X3_Y0                (CDIDATA_X3_Y0_D2),
    .CDIVALID_X3_Y0               (CDIVALID_X3_Y0_D2),
    .CDIREADY_X3_Y0               (CDIREADY_X3_Y0_D2),
    .CDODATA_X3_Y0                (CDODATA_X3_Y0_D2),
    .CDOVALID_X3_Y0               (CDOVALID_X3_Y0_D2),
    .CDOREADY_X3_Y0               (CDOREADY_X3_Y0_D2),
    .CDIDATA_X3_Y1                (CDIDATA_X3_Y1_D2),
    .CDIVALID_X3_Y1               (CDIVALID_X3_Y1_D2),
    .CDIREADY_X3_Y1               (CDIREADY_X3_Y1_D2),
    .CDODATA_X3_Y1                (CDODATA_X3_Y1_D2),
    .CDOVALID_X3_Y1               (CDOVALID_X3_Y1_D2),
    .CDOREADY_X3_Y1               (CDOREADY_X3_Y1_D2),
    .CDIDATA_X3_Y2                (CDIDATA_X3_Y2_D2),
    .CDIVALID_X3_Y2               (CDIVALID_X3_Y2_D2),
    .CDIREADY_X3_Y2               (CDIREADY_X3_Y2_D2),
    .CDODATA_X3_Y2                (CDODATA_X3_Y2_D2),
    .CDOVALID_X3_Y2               (CDOVALID_X3_Y2_D2),
    .CDOREADY_X3_Y2               (CDOREADY_X3_Y2_D2),
    .CDIDATA_X3_Y3                (CDIDATA_X3_Y3_D2),
    .CDIVALID_X3_Y3               (CDIVALID_X3_Y3_D2),
    .CDIREADY_X3_Y3               (CDIREADY_X3_Y3_D2),
    .CDODATA_X3_Y3                (CDODATA_X3_Y3_D2),
    .CDOVALID_X3_Y3               (CDOVALID_X3_Y3_D2),
    .CDOREADY_X3_Y3               (CDOREADY_X3_Y3_D2),
    .CDIDATA_X3_Y4                (CDIDATA_X3_Y4_D2),
    .CDIVALID_X3_Y4               (CDIVALID_X3_Y4_D2),
    .CDIREADY_X3_Y4               (CDIREADY_X3_Y4_D2),
    .CDODATA_X3_Y4                (CDODATA_X3_Y4_D2),
    .CDOVALID_X3_Y4               (CDOVALID_X3_Y4_D2),
    .CDOREADY_X3_Y4               (CDOREADY_X3_Y4_D2),
    .CDIDATA_X4_Y0                (CDIDATA_X4_Y0_D2),
    .CDIVALID_X4_Y0               (CDIVALID_X4_Y0_D2),
    .CDIREADY_X4_Y0               (CDIREADY_X4_Y0_D2),
    .CDODATA_X4_Y0                (CDODATA_X4_Y0_D2),
    .CDOVALID_X4_Y0               (CDOVALID_X4_Y0_D2),
    .CDOREADY_X4_Y0               (CDOREADY_X4_Y0_D2),
    .CDIDATA_X4_Y1                (CDIDATA_X4_Y1_D2),
    .CDIVALID_X4_Y1               (CDIVALID_X4_Y1_D2),
    .CDIREADY_X4_Y1               (CDIREADY_X4_Y1_D2),
    .CDODATA_X4_Y1                (CDODATA_X4_Y1_D2),
    .CDOVALID_X4_Y1               (CDOVALID_X4_Y1_D2),
    .CDOREADY_X4_Y1               (CDOREADY_X4_Y1_D2),
    .CDIDATA_X4_Y2                (CDIDATA_X4_Y2_D2),
    .CDIVALID_X4_Y2               (CDIVALID_X4_Y2_D2),
    .CDIREADY_X4_Y2               (CDIREADY_X4_Y2_D2),
    .CDODATA_X4_Y2                (CDODATA_X4_Y2_D2),
    .CDOVALID_X4_Y2               (CDOVALID_X4_Y2_D2),
    .CDOREADY_X4_Y2               (CDOREADY_X4_Y2_D2),
    .CDIDATA_X4_Y3                (CDIDATA_X4_Y3_D2),
    .CDIVALID_X4_Y3               (CDIVALID_X4_Y3_D2),
    .CDIREADY_X4_Y3               (CDIREADY_X4_Y3_D2),
    .CDODATA_X4_Y3                (CDODATA_X4_Y3_D2),
    .CDOVALID_X4_Y3               (CDOVALID_X4_Y3_D2),
    .CDOREADY_X4_Y3               (CDOREADY_X4_Y3_D2),
    .CDIDATA_X4_Y4                (CDIDATA_X4_Y4_D2),
    .CDIVALID_X4_Y4               (CDIVALID_X4_Y4_D2),
    .CDIREADY_X4_Y4               (CDIREADY_X4_Y4_D2),
    .CDODATA_X4_Y4                (CDODATA_X4_Y4_D2),
    .CDOVALID_X4_Y4               (CDOVALID_X4_Y4_D2),
    .CDOREADY_X4_Y4               (CDOREADY_X4_Y4_D2),
    .CPIDATA_W                    (d1_2_d2_data),
    .CPIVALID_W                   (d1_2_d2_valid),
    .CPIREADY_W                   (d1_2_d2_ready),
    .CPODATA_W                    (d2_2_d1_data),
    .CPOVALID_W                   (d2_2_d1_valid),
    .CPOREADY_W                   (d2_2_d1_ready),
    .CPIDATA_E                    (65'b0),
    .CPIVALID_E                   (1'b0),
    .CPIREADY_E                   (),
    .CPODATA_E                    (),
    .CPOVALID_E                   (),
    .CPOREADY_E                   (1'b0)
);

endmodule